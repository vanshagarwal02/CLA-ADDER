magic
tech scmos
timestamp 1731943659
<< nwell >>
rect -470 -32 -438 94
rect -418 -32 -386 94
rect -366 30 -334 94
rect -314 30 -282 94
rect -269 38 -205 102
rect 1161 94 1193 220
rect 1213 94 1245 220
rect 1265 156 1297 220
rect 1317 156 1349 220
rect 1362 164 1426 228
rect 522 -15 584 12
rect 618 -20 645 42
rect 522 -66 584 -39
rect 150 -206 212 -179
rect 246 -211 273 -149
rect 467 -227 521 -165
rect 150 -257 212 -230
rect -437 -427 -405 -301
rect -385 -427 -353 -301
rect -333 -365 -301 -301
rect -281 -365 -249 -301
rect -236 -357 -172 -293
rect 163 -355 217 -293
rect 529 -297 556 -235
rect 712 -334 739 -132
rect 761 -331 788 -269
rect 225 -425 252 -363
rect 1018 -402 1080 -375
rect 1114 -407 1141 -345
rect 1439 -369 1471 -243
rect 1491 -369 1523 -243
rect 1543 -307 1575 -243
rect 1595 -307 1627 -243
rect 1640 -299 1704 -235
rect 1018 -453 1080 -426
rect -546 -806 -514 -680
rect -494 -806 -462 -680
rect -442 -744 -410 -680
rect -390 -744 -358 -680
rect -345 -736 -281 -672
rect 568 -716 622 -654
rect 101 -842 163 -815
rect 197 -847 224 -785
rect 630 -786 657 -724
rect 967 -823 994 -621
rect 1016 -820 1043 -758
rect 1193 -815 1220 -613
rect 1242 -812 1269 -750
rect 1372 -847 1434 -820
rect 1468 -852 1495 -790
rect 101 -893 163 -866
rect 1372 -898 1434 -871
rect 114 -991 168 -929
rect 491 -961 545 -899
rect 709 -961 763 -899
rect 1750 -924 1782 -798
rect 1802 -924 1834 -798
rect 1854 -862 1886 -798
rect 1906 -862 1938 -798
rect 1951 -854 2015 -790
rect -470 -1159 -438 -1033
rect -418 -1159 -386 -1033
rect -366 -1097 -334 -1033
rect -314 -1097 -282 -1033
rect -269 -1089 -205 -1025
rect 176 -1061 203 -999
rect 553 -1031 580 -969
rect 771 -1031 798 -969
rect 566 -1279 620 -1217
rect 628 -1349 655 -1287
rect -479 -1487 -447 -1361
rect -427 -1487 -395 -1361
rect -375 -1425 -343 -1361
rect -323 -1425 -291 -1361
rect -278 -1417 -214 -1353
rect 110 -1502 172 -1475
rect 206 -1507 233 -1445
rect 110 -1553 172 -1526
rect 567 -1562 621 -1500
rect 803 -1509 857 -1447
rect 1146 -1496 1173 -1294
rect 1195 -1493 1222 -1431
rect 123 -1651 177 -1589
rect 629 -1632 656 -1570
rect 865 -1579 892 -1517
rect 185 -1721 212 -1659
rect 812 -1720 866 -1658
rect -495 -1865 -463 -1739
rect -443 -1865 -411 -1739
rect -391 -1803 -359 -1739
rect -339 -1803 -307 -1739
rect -294 -1795 -230 -1731
rect 563 -1833 617 -1771
rect 874 -1790 901 -1728
rect 1157 -1796 1184 -1594
rect 1306 -1660 1333 -1458
rect 1355 -1657 1382 -1595
rect 1206 -1793 1233 -1731
rect 1488 -1811 1550 -1784
rect 1584 -1816 1611 -1754
rect 625 -1903 652 -1841
rect 1488 -1862 1550 -1835
rect 1901 -1874 1933 -1748
rect 1953 -1874 1985 -1748
rect 2005 -1812 2037 -1748
rect 2057 -1812 2089 -1748
rect 2102 -1804 2166 -1740
rect 551 -2082 605 -2020
rect -479 -2235 -447 -2109
rect -427 -2235 -395 -2109
rect -375 -2173 -343 -2109
rect -323 -2173 -291 -2109
rect -278 -2165 -214 -2101
rect 613 -2152 640 -2090
rect 107 -2377 169 -2350
rect 203 -2382 230 -2320
rect 690 -2392 744 -2330
rect 107 -2428 169 -2401
rect 752 -2462 779 -2400
rect 1025 -2444 1079 -2382
rect 120 -2526 174 -2464
rect 1087 -2514 1114 -2452
rect 1355 -2525 1382 -2323
rect 1404 -2522 1431 -2460
rect -470 -2664 -438 -2538
rect -418 -2664 -386 -2538
rect -366 -2602 -334 -2538
rect -314 -2602 -282 -2538
rect -269 -2594 -205 -2530
rect 182 -2596 209 -2534
rect 2090 -2549 2117 -2347
rect 2139 -2546 2166 -2484
rect 2431 -2555 2463 -2429
rect 2483 -2555 2515 -2429
rect 2535 -2493 2567 -2429
rect 2587 -2493 2619 -2429
rect 2632 -2485 2696 -2421
rect 691 -2675 745 -2613
rect 753 -2745 780 -2683
rect 1026 -2727 1080 -2665
rect 1088 -2797 1115 -2735
rect 687 -2946 741 -2884
rect 1362 -2914 1389 -2712
rect 1411 -2911 1438 -2849
rect 749 -3016 776 -2954
rect 1356 -3129 1410 -3067
rect 1654 -3070 1681 -2868
rect 1703 -3067 1730 -3005
rect 675 -3195 729 -3133
rect 1418 -3199 1445 -3137
rect 737 -3265 764 -3203
rect 1016 -3261 1070 -3199
rect 1078 -3331 1105 -3269
rect 692 -3462 746 -3400
rect 754 -3532 781 -3470
rect 680 -3711 734 -3649
rect 742 -3781 769 -3719
<< ntransistor >>
rect 1377 133 1379 153
rect 1409 133 1411 153
rect 1280 109 1282 129
rect 1332 109 1334 129
rect 1176 62 1178 82
rect 1228 62 1230 82
rect 1280 62 1282 82
rect 1332 62 1334 82
rect -254 7 -252 27
rect -222 7 -220 27
rect -351 -17 -349 3
rect -299 -17 -297 3
rect 492 -3 512 -1
rect 595 -15 597 5
rect -455 -64 -453 -44
rect -403 -64 -401 -44
rect -351 -64 -349 -44
rect -299 -64 -297 -44
rect 595 -48 597 -28
rect 631 -50 633 -30
rect 492 -54 512 -52
rect 120 -194 140 -192
rect 223 -206 225 -186
rect 223 -239 225 -219
rect 259 -241 261 -221
rect 120 -245 140 -243
rect 499 -293 501 -253
rect -221 -388 -219 -368
rect -189 -388 -187 -368
rect 499 -358 501 -318
rect 542 -327 544 -307
rect -318 -412 -316 -392
rect -266 -412 -264 -392
rect 195 -421 197 -381
rect 710 -371 712 -351
rect 743 -371 745 -351
rect 774 -361 776 -341
rect 988 -390 1008 -388
rect 1091 -402 1093 -382
rect 1655 -330 1657 -310
rect 1687 -330 1689 -310
rect 1558 -354 1560 -334
rect 1610 -354 1612 -334
rect -422 -459 -420 -439
rect -370 -459 -368 -439
rect -318 -459 -316 -439
rect -266 -459 -264 -439
rect 195 -486 197 -446
rect 238 -455 240 -435
rect 1091 -435 1093 -415
rect 1454 -401 1456 -381
rect 1506 -401 1508 -381
rect 1558 -401 1560 -381
rect 1610 -401 1612 -381
rect 1127 -437 1129 -417
rect 988 -441 1008 -439
rect -330 -767 -328 -747
rect -298 -767 -296 -747
rect -427 -791 -425 -771
rect -375 -791 -373 -771
rect 600 -782 602 -742
rect -531 -838 -529 -818
rect -479 -838 -477 -818
rect -427 -838 -425 -818
rect -375 -838 -373 -818
rect 71 -830 91 -828
rect 174 -842 176 -822
rect 174 -875 176 -855
rect 600 -847 602 -807
rect 643 -816 645 -796
rect 210 -877 212 -857
rect 965 -860 967 -840
rect 998 -860 1000 -840
rect 1029 -850 1031 -830
rect 1191 -852 1193 -832
rect 1224 -852 1226 -832
rect 1255 -842 1257 -822
rect 1342 -835 1362 -833
rect 1445 -847 1447 -827
rect 71 -881 91 -879
rect 1445 -880 1447 -860
rect 1481 -882 1483 -862
rect 1342 -886 1362 -884
rect 1966 -885 1968 -865
rect 1998 -885 2000 -865
rect 1869 -909 1871 -889
rect 1921 -909 1923 -889
rect 146 -1057 148 -1017
rect 523 -1027 525 -987
rect 1765 -956 1767 -936
rect 1817 -956 1819 -936
rect 1869 -956 1871 -936
rect 1921 -956 1923 -936
rect 741 -1027 743 -987
rect -254 -1120 -252 -1100
rect -222 -1120 -220 -1100
rect 146 -1122 148 -1082
rect 189 -1091 191 -1071
rect 523 -1092 525 -1052
rect 566 -1061 568 -1041
rect 741 -1092 743 -1052
rect 784 -1061 786 -1041
rect -351 -1144 -349 -1124
rect -299 -1144 -297 -1124
rect -455 -1191 -453 -1171
rect -403 -1191 -401 -1171
rect -351 -1191 -349 -1171
rect -299 -1191 -297 -1171
rect 598 -1345 600 -1305
rect 598 -1410 600 -1370
rect 641 -1379 643 -1359
rect -263 -1448 -261 -1428
rect -231 -1448 -229 -1428
rect -360 -1472 -358 -1452
rect -308 -1472 -306 -1452
rect 80 -1490 100 -1488
rect -464 -1519 -462 -1499
rect -412 -1519 -410 -1499
rect -360 -1519 -358 -1499
rect -308 -1519 -306 -1499
rect 183 -1502 185 -1482
rect 183 -1535 185 -1515
rect 219 -1537 221 -1517
rect 80 -1541 100 -1539
rect 599 -1628 601 -1588
rect 835 -1575 837 -1535
rect 1144 -1533 1146 -1513
rect 1177 -1533 1179 -1513
rect 1208 -1523 1210 -1503
rect 835 -1640 837 -1600
rect 878 -1609 880 -1589
rect 155 -1717 157 -1677
rect 599 -1693 601 -1653
rect 642 -1662 644 -1642
rect 155 -1782 157 -1742
rect 198 -1751 200 -1731
rect -279 -1826 -277 -1806
rect -247 -1826 -245 -1806
rect 844 -1786 846 -1746
rect -376 -1850 -374 -1830
rect -324 -1850 -322 -1830
rect -480 -1897 -478 -1877
rect -428 -1897 -426 -1877
rect -376 -1897 -374 -1877
rect -324 -1897 -322 -1877
rect 595 -1899 597 -1859
rect 844 -1851 846 -1811
rect 887 -1820 889 -1800
rect 1304 -1697 1306 -1677
rect 1337 -1697 1339 -1677
rect 1368 -1687 1370 -1667
rect 1458 -1799 1478 -1797
rect 1155 -1833 1157 -1813
rect 1188 -1833 1190 -1813
rect 1219 -1823 1221 -1803
rect 1561 -1811 1563 -1791
rect 1561 -1844 1563 -1824
rect 1597 -1846 1599 -1826
rect 1458 -1850 1478 -1848
rect 2117 -1835 2119 -1815
rect 2149 -1835 2151 -1815
rect 2020 -1859 2022 -1839
rect 2072 -1859 2074 -1839
rect 1916 -1906 1918 -1886
rect 1968 -1906 1970 -1886
rect 2020 -1906 2022 -1886
rect 2072 -1906 2074 -1886
rect 595 -1964 597 -1924
rect 638 -1933 640 -1913
rect 583 -2148 585 -2108
rect -263 -2196 -261 -2176
rect -231 -2196 -229 -2176
rect -360 -2220 -358 -2200
rect -308 -2220 -306 -2200
rect 583 -2213 585 -2173
rect 626 -2182 628 -2162
rect -464 -2267 -462 -2247
rect -412 -2267 -410 -2247
rect -360 -2267 -358 -2247
rect -308 -2267 -306 -2247
rect 77 -2365 97 -2363
rect 180 -2377 182 -2357
rect 180 -2410 182 -2390
rect 216 -2412 218 -2392
rect 77 -2416 97 -2414
rect 722 -2458 724 -2418
rect 722 -2523 724 -2483
rect 765 -2492 767 -2472
rect 1057 -2510 1059 -2470
rect 152 -2592 154 -2552
rect -254 -2625 -252 -2605
rect -222 -2625 -220 -2605
rect 1057 -2575 1059 -2535
rect 1100 -2544 1102 -2524
rect 1353 -2562 1355 -2542
rect 1386 -2562 1388 -2542
rect 1417 -2552 1419 -2532
rect 2647 -2516 2649 -2496
rect 2679 -2516 2681 -2496
rect 2550 -2540 2552 -2520
rect 2602 -2540 2604 -2520
rect 2088 -2586 2090 -2566
rect 2121 -2586 2123 -2566
rect 2152 -2576 2154 -2556
rect 2446 -2587 2448 -2567
rect 2498 -2587 2500 -2567
rect 2550 -2587 2552 -2567
rect 2602 -2587 2604 -2567
rect -351 -2649 -349 -2629
rect -299 -2649 -297 -2629
rect 152 -2657 154 -2617
rect 195 -2626 197 -2606
rect -455 -2696 -453 -2676
rect -403 -2696 -401 -2676
rect -351 -2696 -349 -2676
rect -299 -2696 -297 -2676
rect 723 -2741 725 -2701
rect 723 -2806 725 -2766
rect 766 -2775 768 -2755
rect 1058 -2793 1060 -2753
rect 1058 -2858 1060 -2818
rect 1101 -2827 1103 -2807
rect 1360 -2951 1362 -2931
rect 1393 -2951 1395 -2931
rect 1424 -2941 1426 -2921
rect 719 -3012 721 -2972
rect 719 -3077 721 -3037
rect 762 -3046 764 -3026
rect 1652 -3107 1654 -3087
rect 1685 -3107 1687 -3087
rect 1716 -3097 1718 -3077
rect 1388 -3195 1390 -3155
rect 707 -3261 709 -3221
rect 707 -3326 709 -3286
rect 750 -3295 752 -3275
rect 1388 -3260 1390 -3220
rect 1431 -3229 1433 -3209
rect 1048 -3327 1050 -3287
rect 1048 -3392 1050 -3352
rect 1091 -3361 1093 -3341
rect 724 -3528 726 -3488
rect 724 -3593 726 -3553
rect 767 -3562 769 -3542
rect 712 -3777 714 -3737
rect 712 -3842 714 -3802
rect 755 -3811 757 -3791
<< ptransistor >>
rect 1176 165 1178 205
rect 1228 165 1230 205
rect 1280 165 1282 205
rect 1332 165 1334 205
rect 1377 173 1379 213
rect 1409 173 1411 213
rect 1176 103 1178 143
rect 1228 103 1230 143
rect -455 39 -453 79
rect -403 39 -401 79
rect -351 39 -349 79
rect -299 39 -297 79
rect -254 47 -252 87
rect -222 47 -220 87
rect -455 -23 -453 17
rect -403 -23 -401 17
rect 530 -3 570 -1
rect 631 -12 633 28
rect 530 -54 570 -52
rect 158 -194 198 -192
rect 259 -203 261 -163
rect 480 -219 482 -179
rect 507 -219 509 -179
rect 158 -245 198 -243
rect 725 -226 727 -146
rect -422 -356 -420 -316
rect -370 -356 -368 -316
rect -318 -356 -316 -316
rect -266 -356 -264 -316
rect -221 -348 -219 -308
rect -189 -348 -187 -308
rect 176 -347 178 -307
rect 203 -347 205 -307
rect 542 -289 544 -249
rect -422 -418 -420 -378
rect -370 -418 -368 -378
rect 725 -326 727 -246
rect 774 -323 776 -283
rect 1454 -298 1456 -258
rect 1506 -298 1508 -258
rect 1558 -298 1560 -258
rect 1610 -298 1612 -258
rect 1655 -290 1657 -250
rect 1687 -290 1689 -250
rect 238 -417 240 -377
rect 1026 -390 1066 -388
rect 1127 -399 1129 -359
rect 1454 -360 1456 -320
rect 1506 -360 1508 -320
rect 1026 -441 1066 -439
rect -531 -735 -529 -695
rect -479 -735 -477 -695
rect -427 -735 -425 -695
rect -375 -735 -373 -695
rect -330 -727 -328 -687
rect -298 -727 -296 -687
rect 581 -708 583 -668
rect 608 -708 610 -668
rect 980 -715 982 -635
rect 1206 -707 1208 -627
rect -531 -797 -529 -757
rect -479 -797 -477 -757
rect 643 -778 645 -738
rect 109 -830 149 -828
rect 210 -839 212 -799
rect 980 -815 982 -735
rect 1029 -812 1031 -772
rect 1206 -807 1208 -727
rect 1255 -804 1257 -764
rect 1380 -835 1420 -833
rect 1481 -844 1483 -804
rect 109 -881 149 -879
rect 1765 -853 1767 -813
rect 1817 -853 1819 -813
rect 1869 -853 1871 -813
rect 1921 -853 1923 -813
rect 1966 -845 1968 -805
rect 1998 -845 2000 -805
rect 1380 -886 1420 -884
rect 127 -983 129 -943
rect 154 -983 156 -943
rect 504 -953 506 -913
rect 531 -953 533 -913
rect 722 -953 724 -913
rect 749 -953 751 -913
rect 1765 -915 1767 -875
rect 1817 -915 1819 -875
rect -455 -1088 -453 -1048
rect -403 -1088 -401 -1048
rect -351 -1088 -349 -1048
rect -299 -1088 -297 -1048
rect -254 -1080 -252 -1040
rect -222 -1080 -220 -1040
rect 189 -1053 191 -1013
rect 566 -1023 568 -983
rect -455 -1150 -453 -1110
rect -403 -1150 -401 -1110
rect 784 -1023 786 -983
rect 579 -1271 581 -1231
rect 606 -1271 608 -1231
rect 641 -1341 643 -1301
rect -464 -1416 -462 -1376
rect -412 -1416 -410 -1376
rect -360 -1416 -358 -1376
rect -308 -1416 -306 -1376
rect -263 -1408 -261 -1368
rect -231 -1408 -229 -1368
rect 1159 -1388 1161 -1308
rect -464 -1478 -462 -1438
rect -412 -1478 -410 -1438
rect 118 -1490 158 -1488
rect 219 -1499 221 -1459
rect 816 -1501 818 -1461
rect 843 -1501 845 -1461
rect 1159 -1488 1161 -1408
rect 118 -1541 158 -1539
rect 580 -1554 582 -1514
rect 607 -1554 609 -1514
rect 1208 -1485 1210 -1445
rect 136 -1643 138 -1603
rect 163 -1643 165 -1603
rect 642 -1624 644 -1584
rect 878 -1571 880 -1531
rect 1319 -1552 1321 -1472
rect 198 -1713 200 -1673
rect 825 -1712 827 -1672
rect 852 -1712 854 -1672
rect 1170 -1688 1172 -1608
rect 1319 -1652 1321 -1572
rect 1368 -1649 1370 -1609
rect -480 -1794 -478 -1754
rect -428 -1794 -426 -1754
rect -376 -1794 -374 -1754
rect -324 -1794 -322 -1754
rect -279 -1786 -277 -1746
rect -247 -1786 -245 -1746
rect -480 -1856 -478 -1816
rect -428 -1856 -426 -1816
rect 576 -1825 578 -1785
rect 603 -1825 605 -1785
rect 887 -1782 889 -1742
rect 1170 -1788 1172 -1708
rect 1219 -1785 1221 -1745
rect 1496 -1799 1536 -1797
rect 1597 -1808 1599 -1768
rect 1916 -1803 1918 -1763
rect 1968 -1803 1970 -1763
rect 2020 -1803 2022 -1763
rect 2072 -1803 2074 -1763
rect 2117 -1795 2119 -1755
rect 2149 -1795 2151 -1755
rect 1496 -1850 1536 -1848
rect 638 -1895 640 -1855
rect 1916 -1865 1918 -1825
rect 1968 -1865 1970 -1825
rect 564 -2074 566 -2034
rect 591 -2074 593 -2034
rect -464 -2164 -462 -2124
rect -412 -2164 -410 -2124
rect -360 -2164 -358 -2124
rect -308 -2164 -306 -2124
rect -263 -2156 -261 -2116
rect -231 -2156 -229 -2116
rect 626 -2144 628 -2104
rect -464 -2226 -462 -2186
rect -412 -2226 -410 -2186
rect 115 -2365 155 -2363
rect 216 -2374 218 -2334
rect 703 -2384 705 -2344
rect 730 -2384 732 -2344
rect 115 -2416 155 -2414
rect 765 -2454 767 -2414
rect 1038 -2436 1040 -2396
rect 1065 -2436 1067 -2396
rect 1368 -2417 1370 -2337
rect 133 -2518 135 -2478
rect 160 -2518 162 -2478
rect -455 -2593 -453 -2553
rect -403 -2593 -401 -2553
rect -351 -2593 -349 -2553
rect -299 -2593 -297 -2553
rect -254 -2585 -252 -2545
rect -222 -2585 -220 -2545
rect 1100 -2506 1102 -2466
rect 1368 -2517 1370 -2437
rect -455 -2655 -453 -2615
rect -403 -2655 -401 -2615
rect 195 -2588 197 -2548
rect 2103 -2441 2105 -2361
rect 1417 -2514 1419 -2474
rect 2103 -2541 2105 -2461
rect 2446 -2484 2448 -2444
rect 2498 -2484 2500 -2444
rect 2550 -2484 2552 -2444
rect 2602 -2484 2604 -2444
rect 2647 -2476 2649 -2436
rect 2679 -2476 2681 -2436
rect 2152 -2538 2154 -2498
rect 2446 -2546 2448 -2506
rect 2498 -2546 2500 -2506
rect 704 -2667 706 -2627
rect 731 -2667 733 -2627
rect 766 -2737 768 -2697
rect 1039 -2719 1041 -2679
rect 1066 -2719 1068 -2679
rect 1101 -2789 1103 -2749
rect 1375 -2806 1377 -2726
rect 700 -2938 702 -2898
rect 727 -2938 729 -2898
rect 1375 -2906 1377 -2826
rect 1424 -2903 1426 -2863
rect 1667 -2962 1669 -2882
rect 762 -3008 764 -2968
rect 1667 -3062 1669 -2982
rect 1369 -3121 1371 -3081
rect 1396 -3121 1398 -3081
rect 1716 -3059 1718 -3019
rect 688 -3187 690 -3147
rect 715 -3187 717 -3147
rect 1431 -3191 1433 -3151
rect 750 -3257 752 -3217
rect 1029 -3253 1031 -3213
rect 1056 -3253 1058 -3213
rect 1091 -3323 1093 -3283
rect 705 -3454 707 -3414
rect 732 -3454 734 -3414
rect 767 -3524 769 -3484
rect 693 -3703 695 -3663
rect 720 -3703 722 -3663
rect 755 -3773 757 -3733
<< ndiffusion >>
rect 1376 133 1377 153
rect 1379 133 1380 153
rect 1408 133 1409 153
rect 1411 133 1412 153
rect 1279 109 1280 129
rect 1282 109 1283 129
rect 1331 109 1332 129
rect 1334 109 1335 129
rect 1175 62 1176 82
rect 1178 62 1179 82
rect 1227 62 1228 82
rect 1230 62 1231 82
rect 1279 62 1280 82
rect 1282 62 1283 82
rect 1331 62 1332 82
rect 1334 62 1335 82
rect -255 7 -254 27
rect -252 7 -251 27
rect -223 7 -222 27
rect -220 7 -219 27
rect -352 -17 -351 3
rect -349 -17 -348 3
rect -300 -17 -299 3
rect -297 -17 -296 3
rect 492 -1 512 0
rect 492 -4 512 -3
rect 594 -15 595 5
rect 597 -15 598 5
rect -456 -64 -455 -44
rect -453 -64 -452 -44
rect -404 -64 -403 -44
rect -401 -64 -400 -44
rect -352 -64 -351 -44
rect -349 -64 -348 -44
rect -300 -64 -299 -44
rect -297 -64 -296 -44
rect 492 -52 512 -51
rect 594 -48 595 -28
rect 597 -48 598 -28
rect 630 -50 631 -30
rect 633 -50 634 -30
rect 492 -55 512 -54
rect 120 -192 140 -191
rect 120 -195 140 -194
rect 222 -206 223 -186
rect 225 -206 226 -186
rect 120 -243 140 -242
rect 222 -239 223 -219
rect 225 -239 226 -219
rect 258 -241 259 -221
rect 261 -241 262 -221
rect 120 -246 140 -245
rect 498 -293 499 -253
rect 501 -293 502 -253
rect -222 -388 -221 -368
rect -219 -388 -218 -368
rect -190 -388 -189 -368
rect -187 -388 -186 -368
rect 498 -358 499 -318
rect 501 -358 502 -318
rect 541 -327 542 -307
rect 544 -327 545 -307
rect -319 -412 -318 -392
rect -316 -412 -315 -392
rect -267 -412 -266 -392
rect -264 -412 -263 -392
rect 194 -421 195 -381
rect 197 -421 198 -381
rect 709 -371 710 -351
rect 712 -371 713 -351
rect 742 -371 743 -351
rect 745 -371 746 -351
rect 773 -361 774 -341
rect 776 -361 777 -341
rect 988 -388 1008 -387
rect 988 -391 1008 -390
rect 1090 -402 1091 -382
rect 1093 -402 1094 -382
rect 1654 -330 1655 -310
rect 1657 -330 1658 -310
rect 1686 -330 1687 -310
rect 1689 -330 1690 -310
rect 1557 -354 1558 -334
rect 1560 -354 1561 -334
rect 1609 -354 1610 -334
rect 1612 -354 1613 -334
rect -423 -459 -422 -439
rect -420 -459 -419 -439
rect -371 -459 -370 -439
rect -368 -459 -367 -439
rect -319 -459 -318 -439
rect -316 -459 -315 -439
rect -267 -459 -266 -439
rect -264 -459 -263 -439
rect 194 -486 195 -446
rect 197 -486 198 -446
rect 237 -455 238 -435
rect 240 -455 241 -435
rect 988 -439 1008 -438
rect 1090 -435 1091 -415
rect 1093 -435 1094 -415
rect 1453 -401 1454 -381
rect 1456 -401 1457 -381
rect 1505 -401 1506 -381
rect 1508 -401 1509 -381
rect 1557 -401 1558 -381
rect 1560 -401 1561 -381
rect 1609 -401 1610 -381
rect 1612 -401 1613 -381
rect 1126 -437 1127 -417
rect 1129 -437 1130 -417
rect 988 -442 1008 -441
rect -331 -767 -330 -747
rect -328 -767 -327 -747
rect -299 -767 -298 -747
rect -296 -767 -295 -747
rect -428 -791 -427 -771
rect -425 -791 -424 -771
rect -376 -791 -375 -771
rect -373 -791 -372 -771
rect 599 -782 600 -742
rect 602 -782 603 -742
rect -532 -838 -531 -818
rect -529 -838 -528 -818
rect -480 -838 -479 -818
rect -477 -838 -476 -818
rect -428 -838 -427 -818
rect -425 -838 -424 -818
rect -376 -838 -375 -818
rect -373 -838 -372 -818
rect 71 -828 91 -827
rect 71 -831 91 -830
rect 173 -842 174 -822
rect 176 -842 177 -822
rect 71 -879 91 -878
rect 173 -875 174 -855
rect 176 -875 177 -855
rect 599 -847 600 -807
rect 602 -847 603 -807
rect 642 -816 643 -796
rect 645 -816 646 -796
rect 209 -877 210 -857
rect 212 -877 213 -857
rect 964 -860 965 -840
rect 967 -860 968 -840
rect 997 -860 998 -840
rect 1000 -860 1001 -840
rect 1028 -850 1029 -830
rect 1031 -850 1032 -830
rect 1190 -852 1191 -832
rect 1193 -852 1194 -832
rect 1223 -852 1224 -832
rect 1226 -852 1227 -832
rect 1254 -842 1255 -822
rect 1257 -842 1258 -822
rect 1342 -833 1362 -832
rect 1342 -836 1362 -835
rect 1444 -847 1445 -827
rect 1447 -847 1448 -827
rect 71 -882 91 -881
rect 1342 -884 1362 -883
rect 1444 -880 1445 -860
rect 1447 -880 1448 -860
rect 1480 -882 1481 -862
rect 1483 -882 1484 -862
rect 1342 -887 1362 -886
rect 1965 -885 1966 -865
rect 1968 -885 1969 -865
rect 1997 -885 1998 -865
rect 2000 -885 2001 -865
rect 1868 -909 1869 -889
rect 1871 -909 1872 -889
rect 1920 -909 1921 -889
rect 1923 -909 1924 -889
rect 145 -1057 146 -1017
rect 148 -1057 149 -1017
rect 522 -1027 523 -987
rect 525 -1027 526 -987
rect 1764 -956 1765 -936
rect 1767 -956 1768 -936
rect 1816 -956 1817 -936
rect 1819 -956 1820 -936
rect 1868 -956 1869 -936
rect 1871 -956 1872 -936
rect 1920 -956 1921 -936
rect 1923 -956 1924 -936
rect 740 -1027 741 -987
rect 743 -1027 744 -987
rect -255 -1120 -254 -1100
rect -252 -1120 -251 -1100
rect -223 -1120 -222 -1100
rect -220 -1120 -219 -1100
rect 145 -1122 146 -1082
rect 148 -1122 149 -1082
rect 188 -1091 189 -1071
rect 191 -1091 192 -1071
rect 522 -1092 523 -1052
rect 525 -1092 526 -1052
rect 565 -1061 566 -1041
rect 568 -1061 569 -1041
rect 740 -1092 741 -1052
rect 743 -1092 744 -1052
rect 783 -1061 784 -1041
rect 786 -1061 787 -1041
rect -352 -1144 -351 -1124
rect -349 -1144 -348 -1124
rect -300 -1144 -299 -1124
rect -297 -1144 -296 -1124
rect -456 -1191 -455 -1171
rect -453 -1191 -452 -1171
rect -404 -1191 -403 -1171
rect -401 -1191 -400 -1171
rect -352 -1191 -351 -1171
rect -349 -1191 -348 -1171
rect -300 -1191 -299 -1171
rect -297 -1191 -296 -1171
rect 597 -1345 598 -1305
rect 600 -1345 601 -1305
rect 597 -1410 598 -1370
rect 600 -1410 601 -1370
rect 640 -1379 641 -1359
rect 643 -1379 644 -1359
rect -264 -1448 -263 -1428
rect -261 -1448 -260 -1428
rect -232 -1448 -231 -1428
rect -229 -1448 -228 -1428
rect -361 -1472 -360 -1452
rect -358 -1472 -357 -1452
rect -309 -1472 -308 -1452
rect -306 -1472 -305 -1452
rect 80 -1488 100 -1487
rect 80 -1491 100 -1490
rect -465 -1519 -464 -1499
rect -462 -1519 -461 -1499
rect -413 -1519 -412 -1499
rect -410 -1519 -409 -1499
rect -361 -1519 -360 -1499
rect -358 -1519 -357 -1499
rect -309 -1519 -308 -1499
rect -306 -1519 -305 -1499
rect 182 -1502 183 -1482
rect 185 -1502 186 -1482
rect 80 -1539 100 -1538
rect 182 -1535 183 -1515
rect 185 -1535 186 -1515
rect 218 -1537 219 -1517
rect 221 -1537 222 -1517
rect 80 -1542 100 -1541
rect 598 -1628 599 -1588
rect 601 -1628 602 -1588
rect 834 -1575 835 -1535
rect 837 -1575 838 -1535
rect 1143 -1533 1144 -1513
rect 1146 -1533 1147 -1513
rect 1176 -1533 1177 -1513
rect 1179 -1533 1180 -1513
rect 1207 -1523 1208 -1503
rect 1210 -1523 1211 -1503
rect 834 -1640 835 -1600
rect 837 -1640 838 -1600
rect 877 -1609 878 -1589
rect 880 -1609 881 -1589
rect 154 -1717 155 -1677
rect 157 -1717 158 -1677
rect 598 -1693 599 -1653
rect 601 -1693 602 -1653
rect 641 -1662 642 -1642
rect 644 -1662 645 -1642
rect 154 -1782 155 -1742
rect 157 -1782 158 -1742
rect 197 -1751 198 -1731
rect 200 -1751 201 -1731
rect -280 -1826 -279 -1806
rect -277 -1826 -276 -1806
rect -248 -1826 -247 -1806
rect -245 -1826 -244 -1806
rect 843 -1786 844 -1746
rect 846 -1786 847 -1746
rect -377 -1850 -376 -1830
rect -374 -1850 -373 -1830
rect -325 -1850 -324 -1830
rect -322 -1850 -321 -1830
rect -481 -1897 -480 -1877
rect -478 -1897 -477 -1877
rect -429 -1897 -428 -1877
rect -426 -1897 -425 -1877
rect -377 -1897 -376 -1877
rect -374 -1897 -373 -1877
rect -325 -1897 -324 -1877
rect -322 -1897 -321 -1877
rect 594 -1899 595 -1859
rect 597 -1899 598 -1859
rect 843 -1851 844 -1811
rect 846 -1851 847 -1811
rect 886 -1820 887 -1800
rect 889 -1820 890 -1800
rect 1303 -1697 1304 -1677
rect 1306 -1697 1307 -1677
rect 1336 -1697 1337 -1677
rect 1339 -1697 1340 -1677
rect 1367 -1687 1368 -1667
rect 1370 -1687 1371 -1667
rect 1458 -1797 1478 -1796
rect 1458 -1800 1478 -1799
rect 1154 -1833 1155 -1813
rect 1157 -1833 1158 -1813
rect 1187 -1833 1188 -1813
rect 1190 -1833 1191 -1813
rect 1218 -1823 1219 -1803
rect 1221 -1823 1222 -1803
rect 1560 -1811 1561 -1791
rect 1563 -1811 1564 -1791
rect 1458 -1848 1478 -1847
rect 1560 -1844 1561 -1824
rect 1563 -1844 1564 -1824
rect 1596 -1846 1597 -1826
rect 1599 -1846 1600 -1826
rect 1458 -1851 1478 -1850
rect 2116 -1835 2117 -1815
rect 2119 -1835 2120 -1815
rect 2148 -1835 2149 -1815
rect 2151 -1835 2152 -1815
rect 2019 -1859 2020 -1839
rect 2022 -1859 2023 -1839
rect 2071 -1859 2072 -1839
rect 2074 -1859 2075 -1839
rect 1915 -1906 1916 -1886
rect 1918 -1906 1919 -1886
rect 1967 -1906 1968 -1886
rect 1970 -1906 1971 -1886
rect 2019 -1906 2020 -1886
rect 2022 -1906 2023 -1886
rect 2071 -1906 2072 -1886
rect 2074 -1906 2075 -1886
rect 594 -1964 595 -1924
rect 597 -1964 598 -1924
rect 637 -1933 638 -1913
rect 640 -1933 641 -1913
rect 582 -2148 583 -2108
rect 585 -2148 586 -2108
rect -264 -2196 -263 -2176
rect -261 -2196 -260 -2176
rect -232 -2196 -231 -2176
rect -229 -2196 -228 -2176
rect -361 -2220 -360 -2200
rect -358 -2220 -357 -2200
rect -309 -2220 -308 -2200
rect -306 -2220 -305 -2200
rect 582 -2213 583 -2173
rect 585 -2213 586 -2173
rect 625 -2182 626 -2162
rect 628 -2182 629 -2162
rect -465 -2267 -464 -2247
rect -462 -2267 -461 -2247
rect -413 -2267 -412 -2247
rect -410 -2267 -409 -2247
rect -361 -2267 -360 -2247
rect -358 -2267 -357 -2247
rect -309 -2267 -308 -2247
rect -306 -2267 -305 -2247
rect 77 -2363 97 -2362
rect 77 -2366 97 -2365
rect 179 -2377 180 -2357
rect 182 -2377 183 -2357
rect 77 -2414 97 -2413
rect 179 -2410 180 -2390
rect 182 -2410 183 -2390
rect 215 -2412 216 -2392
rect 218 -2412 219 -2392
rect 77 -2417 97 -2416
rect 721 -2458 722 -2418
rect 724 -2458 725 -2418
rect 721 -2523 722 -2483
rect 724 -2523 725 -2483
rect 764 -2492 765 -2472
rect 767 -2492 768 -2472
rect 1056 -2510 1057 -2470
rect 1059 -2510 1060 -2470
rect 151 -2592 152 -2552
rect 154 -2592 155 -2552
rect -255 -2625 -254 -2605
rect -252 -2625 -251 -2605
rect -223 -2625 -222 -2605
rect -220 -2625 -219 -2605
rect 1056 -2575 1057 -2535
rect 1059 -2575 1060 -2535
rect 1099 -2544 1100 -2524
rect 1102 -2544 1103 -2524
rect 1352 -2562 1353 -2542
rect 1355 -2562 1356 -2542
rect 1385 -2562 1386 -2542
rect 1388 -2562 1389 -2542
rect 1416 -2552 1417 -2532
rect 1419 -2552 1420 -2532
rect 2646 -2516 2647 -2496
rect 2649 -2516 2650 -2496
rect 2678 -2516 2679 -2496
rect 2681 -2516 2682 -2496
rect 2549 -2540 2550 -2520
rect 2552 -2540 2553 -2520
rect 2601 -2540 2602 -2520
rect 2604 -2540 2605 -2520
rect 2087 -2586 2088 -2566
rect 2090 -2586 2091 -2566
rect 2120 -2586 2121 -2566
rect 2123 -2586 2124 -2566
rect 2151 -2576 2152 -2556
rect 2154 -2576 2155 -2556
rect 2445 -2587 2446 -2567
rect 2448 -2587 2449 -2567
rect 2497 -2587 2498 -2567
rect 2500 -2587 2501 -2567
rect 2549 -2587 2550 -2567
rect 2552 -2587 2553 -2567
rect 2601 -2587 2602 -2567
rect 2604 -2587 2605 -2567
rect -352 -2649 -351 -2629
rect -349 -2649 -348 -2629
rect -300 -2649 -299 -2629
rect -297 -2649 -296 -2629
rect 151 -2657 152 -2617
rect 154 -2657 155 -2617
rect 194 -2626 195 -2606
rect 197 -2626 198 -2606
rect -456 -2696 -455 -2676
rect -453 -2696 -452 -2676
rect -404 -2696 -403 -2676
rect -401 -2696 -400 -2676
rect -352 -2696 -351 -2676
rect -349 -2696 -348 -2676
rect -300 -2696 -299 -2676
rect -297 -2696 -296 -2676
rect 722 -2741 723 -2701
rect 725 -2741 726 -2701
rect 722 -2806 723 -2766
rect 725 -2806 726 -2766
rect 765 -2775 766 -2755
rect 768 -2775 769 -2755
rect 1057 -2793 1058 -2753
rect 1060 -2793 1061 -2753
rect 1057 -2858 1058 -2818
rect 1060 -2858 1061 -2818
rect 1100 -2827 1101 -2807
rect 1103 -2827 1104 -2807
rect 1359 -2951 1360 -2931
rect 1362 -2951 1363 -2931
rect 1392 -2951 1393 -2931
rect 1395 -2951 1396 -2931
rect 1423 -2941 1424 -2921
rect 1426 -2941 1427 -2921
rect 718 -3012 719 -2972
rect 721 -3012 722 -2972
rect 718 -3077 719 -3037
rect 721 -3077 722 -3037
rect 761 -3046 762 -3026
rect 764 -3046 765 -3026
rect 1651 -3107 1652 -3087
rect 1654 -3107 1655 -3087
rect 1684 -3107 1685 -3087
rect 1687 -3107 1688 -3087
rect 1715 -3097 1716 -3077
rect 1718 -3097 1719 -3077
rect 1387 -3195 1388 -3155
rect 1390 -3195 1391 -3155
rect 706 -3261 707 -3221
rect 709 -3261 710 -3221
rect 706 -3326 707 -3286
rect 709 -3326 710 -3286
rect 749 -3295 750 -3275
rect 752 -3295 753 -3275
rect 1387 -3260 1388 -3220
rect 1390 -3260 1391 -3220
rect 1430 -3229 1431 -3209
rect 1433 -3229 1434 -3209
rect 1047 -3327 1048 -3287
rect 1050 -3327 1051 -3287
rect 1047 -3392 1048 -3352
rect 1050 -3392 1051 -3352
rect 1090 -3361 1091 -3341
rect 1093 -3361 1094 -3341
rect 723 -3528 724 -3488
rect 726 -3528 727 -3488
rect 723 -3593 724 -3553
rect 726 -3593 727 -3553
rect 766 -3562 767 -3542
rect 769 -3562 770 -3542
rect 711 -3777 712 -3737
rect 714 -3777 715 -3737
rect 711 -3842 712 -3802
rect 714 -3842 715 -3802
rect 754 -3811 755 -3791
rect 757 -3811 758 -3791
<< pdiffusion >>
rect 1175 165 1176 205
rect 1178 165 1179 205
rect 1227 165 1228 205
rect 1230 165 1231 205
rect 1279 165 1280 205
rect 1282 165 1283 205
rect 1331 165 1332 205
rect 1334 165 1335 205
rect 1376 173 1377 213
rect 1379 173 1380 213
rect 1408 173 1409 213
rect 1411 173 1412 213
rect 1175 103 1176 143
rect 1178 103 1179 143
rect 1227 103 1228 143
rect 1230 103 1231 143
rect -456 39 -455 79
rect -453 39 -452 79
rect -404 39 -403 79
rect -401 39 -400 79
rect -352 39 -351 79
rect -349 39 -348 79
rect -300 39 -299 79
rect -297 39 -296 79
rect -255 47 -254 87
rect -252 47 -251 87
rect -223 47 -222 87
rect -220 47 -219 87
rect -456 -23 -455 17
rect -453 -23 -452 17
rect -404 -23 -403 17
rect -401 -23 -400 17
rect 530 -1 570 0
rect 530 -4 570 -3
rect 630 -12 631 28
rect 633 -12 634 28
rect 530 -52 570 -51
rect 530 -55 570 -54
rect 158 -192 198 -191
rect 158 -195 198 -194
rect 258 -203 259 -163
rect 261 -203 262 -163
rect 479 -219 480 -179
rect 482 -219 483 -179
rect 506 -219 507 -179
rect 509 -219 510 -179
rect 158 -243 198 -242
rect 158 -246 198 -245
rect 724 -226 725 -146
rect 727 -226 728 -146
rect -423 -356 -422 -316
rect -420 -356 -419 -316
rect -371 -356 -370 -316
rect -368 -356 -367 -316
rect -319 -356 -318 -316
rect -316 -356 -315 -316
rect -267 -356 -266 -316
rect -264 -356 -263 -316
rect -222 -348 -221 -308
rect -219 -348 -218 -308
rect -190 -348 -189 -308
rect -187 -348 -186 -308
rect 175 -347 176 -307
rect 178 -347 179 -307
rect 202 -347 203 -307
rect 205 -347 206 -307
rect 541 -289 542 -249
rect 544 -289 545 -249
rect -423 -418 -422 -378
rect -420 -418 -419 -378
rect -371 -418 -370 -378
rect -368 -418 -367 -378
rect 724 -326 725 -246
rect 727 -326 728 -246
rect 773 -323 774 -283
rect 776 -323 777 -283
rect 1453 -298 1454 -258
rect 1456 -298 1457 -258
rect 1505 -298 1506 -258
rect 1508 -298 1509 -258
rect 1557 -298 1558 -258
rect 1560 -298 1561 -258
rect 1609 -298 1610 -258
rect 1612 -298 1613 -258
rect 1654 -290 1655 -250
rect 1657 -290 1658 -250
rect 1686 -290 1687 -250
rect 1689 -290 1690 -250
rect 237 -417 238 -377
rect 240 -417 241 -377
rect 1026 -388 1066 -387
rect 1026 -391 1066 -390
rect 1126 -399 1127 -359
rect 1129 -399 1130 -359
rect 1453 -360 1454 -320
rect 1456 -360 1457 -320
rect 1505 -360 1506 -320
rect 1508 -360 1509 -320
rect 1026 -439 1066 -438
rect 1026 -442 1066 -441
rect -532 -735 -531 -695
rect -529 -735 -528 -695
rect -480 -735 -479 -695
rect -477 -735 -476 -695
rect -428 -735 -427 -695
rect -425 -735 -424 -695
rect -376 -735 -375 -695
rect -373 -735 -372 -695
rect -331 -727 -330 -687
rect -328 -727 -327 -687
rect -299 -727 -298 -687
rect -296 -727 -295 -687
rect 580 -708 581 -668
rect 583 -708 584 -668
rect 607 -708 608 -668
rect 610 -708 611 -668
rect 979 -715 980 -635
rect 982 -715 983 -635
rect 1205 -707 1206 -627
rect 1208 -707 1209 -627
rect -532 -797 -531 -757
rect -529 -797 -528 -757
rect -480 -797 -479 -757
rect -477 -797 -476 -757
rect 642 -778 643 -738
rect 645 -778 646 -738
rect 109 -828 149 -827
rect 109 -831 149 -830
rect 209 -839 210 -799
rect 212 -839 213 -799
rect 979 -815 980 -735
rect 982 -815 983 -735
rect 1028 -812 1029 -772
rect 1031 -812 1032 -772
rect 1205 -807 1206 -727
rect 1208 -807 1209 -727
rect 1254 -804 1255 -764
rect 1257 -804 1258 -764
rect 1380 -833 1420 -832
rect 1380 -836 1420 -835
rect 1480 -844 1481 -804
rect 1483 -844 1484 -804
rect 109 -879 149 -878
rect 109 -882 149 -881
rect 1764 -853 1765 -813
rect 1767 -853 1768 -813
rect 1816 -853 1817 -813
rect 1819 -853 1820 -813
rect 1868 -853 1869 -813
rect 1871 -853 1872 -813
rect 1920 -853 1921 -813
rect 1923 -853 1924 -813
rect 1965 -845 1966 -805
rect 1968 -845 1969 -805
rect 1997 -845 1998 -805
rect 2000 -845 2001 -805
rect 1380 -884 1420 -883
rect 1380 -887 1420 -886
rect 126 -983 127 -943
rect 129 -983 130 -943
rect 153 -983 154 -943
rect 156 -983 157 -943
rect 503 -953 504 -913
rect 506 -953 507 -913
rect 530 -953 531 -913
rect 533 -953 534 -913
rect 721 -953 722 -913
rect 724 -953 725 -913
rect 748 -953 749 -913
rect 751 -953 752 -913
rect 1764 -915 1765 -875
rect 1767 -915 1768 -875
rect 1816 -915 1817 -875
rect 1819 -915 1820 -875
rect -456 -1088 -455 -1048
rect -453 -1088 -452 -1048
rect -404 -1088 -403 -1048
rect -401 -1088 -400 -1048
rect -352 -1088 -351 -1048
rect -349 -1088 -348 -1048
rect -300 -1088 -299 -1048
rect -297 -1088 -296 -1048
rect -255 -1080 -254 -1040
rect -252 -1080 -251 -1040
rect -223 -1080 -222 -1040
rect -220 -1080 -219 -1040
rect 188 -1053 189 -1013
rect 191 -1053 192 -1013
rect 565 -1023 566 -983
rect 568 -1023 569 -983
rect -456 -1150 -455 -1110
rect -453 -1150 -452 -1110
rect -404 -1150 -403 -1110
rect -401 -1150 -400 -1110
rect 783 -1023 784 -983
rect 786 -1023 787 -983
rect 578 -1271 579 -1231
rect 581 -1271 582 -1231
rect 605 -1271 606 -1231
rect 608 -1271 609 -1231
rect 640 -1341 641 -1301
rect 643 -1341 644 -1301
rect -465 -1416 -464 -1376
rect -462 -1416 -461 -1376
rect -413 -1416 -412 -1376
rect -410 -1416 -409 -1376
rect -361 -1416 -360 -1376
rect -358 -1416 -357 -1376
rect -309 -1416 -308 -1376
rect -306 -1416 -305 -1376
rect -264 -1408 -263 -1368
rect -261 -1408 -260 -1368
rect -232 -1408 -231 -1368
rect -229 -1408 -228 -1368
rect 1158 -1388 1159 -1308
rect 1161 -1388 1162 -1308
rect -465 -1478 -464 -1438
rect -462 -1478 -461 -1438
rect -413 -1478 -412 -1438
rect -410 -1478 -409 -1438
rect 118 -1488 158 -1487
rect 118 -1491 158 -1490
rect 218 -1499 219 -1459
rect 221 -1499 222 -1459
rect 815 -1501 816 -1461
rect 818 -1501 819 -1461
rect 842 -1501 843 -1461
rect 845 -1501 846 -1461
rect 1158 -1488 1159 -1408
rect 1161 -1488 1162 -1408
rect 118 -1539 158 -1538
rect 118 -1542 158 -1541
rect 579 -1554 580 -1514
rect 582 -1554 583 -1514
rect 606 -1554 607 -1514
rect 609 -1554 610 -1514
rect 1207 -1485 1208 -1445
rect 1210 -1485 1211 -1445
rect 135 -1643 136 -1603
rect 138 -1643 139 -1603
rect 162 -1643 163 -1603
rect 165 -1643 166 -1603
rect 641 -1624 642 -1584
rect 644 -1624 645 -1584
rect 877 -1571 878 -1531
rect 880 -1571 881 -1531
rect 1318 -1552 1319 -1472
rect 1321 -1552 1322 -1472
rect 197 -1713 198 -1673
rect 200 -1713 201 -1673
rect 824 -1712 825 -1672
rect 827 -1712 828 -1672
rect 851 -1712 852 -1672
rect 854 -1712 855 -1672
rect 1169 -1688 1170 -1608
rect 1172 -1688 1173 -1608
rect 1318 -1652 1319 -1572
rect 1321 -1652 1322 -1572
rect 1367 -1649 1368 -1609
rect 1370 -1649 1371 -1609
rect -481 -1794 -480 -1754
rect -478 -1794 -477 -1754
rect -429 -1794 -428 -1754
rect -426 -1794 -425 -1754
rect -377 -1794 -376 -1754
rect -374 -1794 -373 -1754
rect -325 -1794 -324 -1754
rect -322 -1794 -321 -1754
rect -280 -1786 -279 -1746
rect -277 -1786 -276 -1746
rect -248 -1786 -247 -1746
rect -245 -1786 -244 -1746
rect -481 -1856 -480 -1816
rect -478 -1856 -477 -1816
rect -429 -1856 -428 -1816
rect -426 -1856 -425 -1816
rect 575 -1825 576 -1785
rect 578 -1825 579 -1785
rect 602 -1825 603 -1785
rect 605 -1825 606 -1785
rect 886 -1782 887 -1742
rect 889 -1782 890 -1742
rect 1169 -1788 1170 -1708
rect 1172 -1788 1173 -1708
rect 1218 -1785 1219 -1745
rect 1221 -1785 1222 -1745
rect 1496 -1797 1536 -1796
rect 1496 -1800 1536 -1799
rect 1596 -1808 1597 -1768
rect 1599 -1808 1600 -1768
rect 1915 -1803 1916 -1763
rect 1918 -1803 1919 -1763
rect 1967 -1803 1968 -1763
rect 1970 -1803 1971 -1763
rect 2019 -1803 2020 -1763
rect 2022 -1803 2023 -1763
rect 2071 -1803 2072 -1763
rect 2074 -1803 2075 -1763
rect 2116 -1795 2117 -1755
rect 2119 -1795 2120 -1755
rect 2148 -1795 2149 -1755
rect 2151 -1795 2152 -1755
rect 1496 -1848 1536 -1847
rect 1496 -1851 1536 -1850
rect 637 -1895 638 -1855
rect 640 -1895 641 -1855
rect 1915 -1865 1916 -1825
rect 1918 -1865 1919 -1825
rect 1967 -1865 1968 -1825
rect 1970 -1865 1971 -1825
rect 563 -2074 564 -2034
rect 566 -2074 567 -2034
rect 590 -2074 591 -2034
rect 593 -2074 594 -2034
rect -465 -2164 -464 -2124
rect -462 -2164 -461 -2124
rect -413 -2164 -412 -2124
rect -410 -2164 -409 -2124
rect -361 -2164 -360 -2124
rect -358 -2164 -357 -2124
rect -309 -2164 -308 -2124
rect -306 -2164 -305 -2124
rect -264 -2156 -263 -2116
rect -261 -2156 -260 -2116
rect -232 -2156 -231 -2116
rect -229 -2156 -228 -2116
rect 625 -2144 626 -2104
rect 628 -2144 629 -2104
rect -465 -2226 -464 -2186
rect -462 -2226 -461 -2186
rect -413 -2226 -412 -2186
rect -410 -2226 -409 -2186
rect 115 -2363 155 -2362
rect 115 -2366 155 -2365
rect 215 -2374 216 -2334
rect 218 -2374 219 -2334
rect 702 -2384 703 -2344
rect 705 -2384 706 -2344
rect 729 -2384 730 -2344
rect 732 -2384 733 -2344
rect 115 -2414 155 -2413
rect 115 -2417 155 -2416
rect 764 -2454 765 -2414
rect 767 -2454 768 -2414
rect 1037 -2436 1038 -2396
rect 1040 -2436 1041 -2396
rect 1064 -2436 1065 -2396
rect 1067 -2436 1068 -2396
rect 1367 -2417 1368 -2337
rect 1370 -2417 1371 -2337
rect 132 -2518 133 -2478
rect 135 -2518 136 -2478
rect 159 -2518 160 -2478
rect 162 -2518 163 -2478
rect -456 -2593 -455 -2553
rect -453 -2593 -452 -2553
rect -404 -2593 -403 -2553
rect -401 -2593 -400 -2553
rect -352 -2593 -351 -2553
rect -349 -2593 -348 -2553
rect -300 -2593 -299 -2553
rect -297 -2593 -296 -2553
rect -255 -2585 -254 -2545
rect -252 -2585 -251 -2545
rect -223 -2585 -222 -2545
rect -220 -2585 -219 -2545
rect 1099 -2506 1100 -2466
rect 1102 -2506 1103 -2466
rect 1367 -2517 1368 -2437
rect 1370 -2517 1371 -2437
rect -456 -2655 -455 -2615
rect -453 -2655 -452 -2615
rect -404 -2655 -403 -2615
rect -401 -2655 -400 -2615
rect 194 -2588 195 -2548
rect 197 -2588 198 -2548
rect 2102 -2441 2103 -2361
rect 2105 -2441 2106 -2361
rect 1416 -2514 1417 -2474
rect 1419 -2514 1420 -2474
rect 2102 -2541 2103 -2461
rect 2105 -2541 2106 -2461
rect 2445 -2484 2446 -2444
rect 2448 -2484 2449 -2444
rect 2497 -2484 2498 -2444
rect 2500 -2484 2501 -2444
rect 2549 -2484 2550 -2444
rect 2552 -2484 2553 -2444
rect 2601 -2484 2602 -2444
rect 2604 -2484 2605 -2444
rect 2646 -2476 2647 -2436
rect 2649 -2476 2650 -2436
rect 2678 -2476 2679 -2436
rect 2681 -2476 2682 -2436
rect 2151 -2538 2152 -2498
rect 2154 -2538 2155 -2498
rect 2445 -2546 2446 -2506
rect 2448 -2546 2449 -2506
rect 2497 -2546 2498 -2506
rect 2500 -2546 2501 -2506
rect 703 -2667 704 -2627
rect 706 -2667 707 -2627
rect 730 -2667 731 -2627
rect 733 -2667 734 -2627
rect 765 -2737 766 -2697
rect 768 -2737 769 -2697
rect 1038 -2719 1039 -2679
rect 1041 -2719 1042 -2679
rect 1065 -2719 1066 -2679
rect 1068 -2719 1069 -2679
rect 1100 -2789 1101 -2749
rect 1103 -2789 1104 -2749
rect 1374 -2806 1375 -2726
rect 1377 -2806 1378 -2726
rect 699 -2938 700 -2898
rect 702 -2938 703 -2898
rect 726 -2938 727 -2898
rect 729 -2938 730 -2898
rect 1374 -2906 1375 -2826
rect 1377 -2906 1378 -2826
rect 1423 -2903 1424 -2863
rect 1426 -2903 1427 -2863
rect 1666 -2962 1667 -2882
rect 1669 -2962 1670 -2882
rect 761 -3008 762 -2968
rect 764 -3008 765 -2968
rect 1666 -3062 1667 -2982
rect 1669 -3062 1670 -2982
rect 1368 -3121 1369 -3081
rect 1371 -3121 1372 -3081
rect 1395 -3121 1396 -3081
rect 1398 -3121 1399 -3081
rect 1715 -3059 1716 -3019
rect 1718 -3059 1719 -3019
rect 687 -3187 688 -3147
rect 690 -3187 691 -3147
rect 714 -3187 715 -3147
rect 717 -3187 718 -3147
rect 1430 -3191 1431 -3151
rect 1433 -3191 1434 -3151
rect 749 -3257 750 -3217
rect 752 -3257 753 -3217
rect 1028 -3253 1029 -3213
rect 1031 -3253 1032 -3213
rect 1055 -3253 1056 -3213
rect 1058 -3253 1059 -3213
rect 1090 -3323 1091 -3283
rect 1093 -3323 1094 -3283
rect 704 -3454 705 -3414
rect 707 -3454 708 -3414
rect 731 -3454 732 -3414
rect 734 -3454 735 -3414
rect 766 -3524 767 -3484
rect 769 -3524 770 -3484
rect 692 -3703 693 -3663
rect 695 -3703 696 -3663
rect 719 -3703 720 -3663
rect 722 -3703 723 -3663
rect 754 -3773 755 -3733
rect 757 -3773 758 -3733
<< ndcontact >>
rect 1372 133 1376 153
rect 1380 133 1384 153
rect 1404 133 1408 153
rect 1412 133 1416 153
rect 1275 109 1279 129
rect 1283 109 1287 129
rect 1327 109 1331 129
rect 1335 109 1339 129
rect 1171 62 1175 82
rect 1179 62 1183 82
rect 1223 62 1227 82
rect 1231 62 1235 82
rect 1275 62 1279 82
rect 1283 62 1287 82
rect 1327 62 1331 82
rect 1335 62 1339 82
rect -259 7 -255 27
rect -251 7 -247 27
rect -227 7 -223 27
rect -219 7 -215 27
rect -356 -17 -352 3
rect -348 -17 -344 3
rect -304 -17 -300 3
rect -296 -17 -292 3
rect 492 0 512 4
rect 492 -8 512 -4
rect 590 -15 594 5
rect 598 -15 602 5
rect -460 -64 -456 -44
rect -452 -64 -448 -44
rect -408 -64 -404 -44
rect -400 -64 -396 -44
rect -356 -64 -352 -44
rect -348 -64 -344 -44
rect -304 -64 -300 -44
rect -296 -64 -292 -44
rect 492 -51 512 -47
rect 590 -48 594 -28
rect 598 -48 602 -28
rect 626 -50 630 -30
rect 634 -50 638 -30
rect 492 -59 512 -55
rect 120 -191 140 -187
rect 120 -199 140 -195
rect 218 -206 222 -186
rect 226 -206 230 -186
rect 120 -242 140 -238
rect 218 -239 222 -219
rect 226 -239 230 -219
rect 254 -241 258 -221
rect 262 -241 266 -221
rect 120 -250 140 -246
rect 494 -293 498 -253
rect 502 -293 506 -253
rect -226 -388 -222 -368
rect -218 -388 -214 -368
rect -194 -388 -190 -368
rect -186 -388 -182 -368
rect 494 -358 498 -318
rect 502 -358 506 -318
rect 537 -327 541 -307
rect 545 -327 549 -307
rect -323 -412 -319 -392
rect -315 -412 -311 -392
rect -271 -412 -267 -392
rect -263 -412 -259 -392
rect 190 -421 194 -381
rect 198 -421 202 -381
rect 705 -371 709 -351
rect 713 -371 717 -351
rect 738 -371 742 -351
rect 746 -371 750 -351
rect 769 -361 773 -341
rect 777 -361 781 -341
rect 988 -387 1008 -383
rect 988 -395 1008 -391
rect 1086 -402 1090 -382
rect 1094 -402 1098 -382
rect 1650 -330 1654 -310
rect 1658 -330 1662 -310
rect 1682 -330 1686 -310
rect 1690 -330 1694 -310
rect 1553 -354 1557 -334
rect 1561 -354 1565 -334
rect 1605 -354 1609 -334
rect 1613 -354 1617 -334
rect -427 -459 -423 -439
rect -419 -459 -415 -439
rect -375 -459 -371 -439
rect -367 -459 -363 -439
rect -323 -459 -319 -439
rect -315 -459 -311 -439
rect -271 -459 -267 -439
rect -263 -459 -259 -439
rect 190 -486 194 -446
rect 198 -486 202 -446
rect 233 -455 237 -435
rect 241 -455 245 -435
rect 988 -438 1008 -434
rect 1086 -435 1090 -415
rect 1094 -435 1098 -415
rect 1449 -401 1453 -381
rect 1457 -401 1461 -381
rect 1501 -401 1505 -381
rect 1509 -401 1513 -381
rect 1553 -401 1557 -381
rect 1561 -401 1565 -381
rect 1605 -401 1609 -381
rect 1613 -401 1617 -381
rect 1122 -437 1126 -417
rect 1130 -437 1134 -417
rect 988 -446 1008 -442
rect -335 -767 -331 -747
rect -327 -767 -323 -747
rect -303 -767 -299 -747
rect -295 -767 -291 -747
rect -432 -791 -428 -771
rect -424 -791 -420 -771
rect -380 -791 -376 -771
rect -372 -791 -368 -771
rect 595 -782 599 -742
rect 603 -782 607 -742
rect -536 -838 -532 -818
rect -528 -838 -524 -818
rect -484 -838 -480 -818
rect -476 -838 -472 -818
rect -432 -838 -428 -818
rect -424 -838 -420 -818
rect -380 -838 -376 -818
rect -372 -838 -368 -818
rect 71 -827 91 -823
rect 71 -835 91 -831
rect 169 -842 173 -822
rect 177 -842 181 -822
rect 71 -878 91 -874
rect 169 -875 173 -855
rect 177 -875 181 -855
rect 595 -847 599 -807
rect 603 -847 607 -807
rect 638 -816 642 -796
rect 646 -816 650 -796
rect 205 -877 209 -857
rect 213 -877 217 -857
rect 960 -860 964 -840
rect 968 -860 972 -840
rect 993 -860 997 -840
rect 1001 -860 1005 -840
rect 1024 -850 1028 -830
rect 1032 -850 1036 -830
rect 1186 -852 1190 -832
rect 1194 -852 1198 -832
rect 1219 -852 1223 -832
rect 1227 -852 1231 -832
rect 1250 -842 1254 -822
rect 1258 -842 1262 -822
rect 1342 -832 1362 -828
rect 1342 -840 1362 -836
rect 1440 -847 1444 -827
rect 1448 -847 1452 -827
rect 71 -886 91 -882
rect 1342 -883 1362 -879
rect 1440 -880 1444 -860
rect 1448 -880 1452 -860
rect 1476 -882 1480 -862
rect 1484 -882 1488 -862
rect 1342 -891 1362 -887
rect 1961 -885 1965 -865
rect 1969 -885 1973 -865
rect 1993 -885 1997 -865
rect 2001 -885 2005 -865
rect 1864 -909 1868 -889
rect 1872 -909 1876 -889
rect 1916 -909 1920 -889
rect 1924 -909 1928 -889
rect 141 -1057 145 -1017
rect 149 -1057 153 -1017
rect 518 -1027 522 -987
rect 526 -1027 530 -987
rect 1760 -956 1764 -936
rect 1768 -956 1772 -936
rect 1812 -956 1816 -936
rect 1820 -956 1824 -936
rect 1864 -956 1868 -936
rect 1872 -956 1876 -936
rect 1916 -956 1920 -936
rect 1924 -956 1928 -936
rect 736 -1027 740 -987
rect 744 -1027 748 -987
rect -259 -1120 -255 -1100
rect -251 -1120 -247 -1100
rect -227 -1120 -223 -1100
rect -219 -1120 -215 -1100
rect 141 -1122 145 -1082
rect 149 -1122 153 -1082
rect 184 -1091 188 -1071
rect 192 -1091 196 -1071
rect 518 -1092 522 -1052
rect 526 -1092 530 -1052
rect 561 -1061 565 -1041
rect 569 -1061 573 -1041
rect 736 -1092 740 -1052
rect 744 -1092 748 -1052
rect 779 -1061 783 -1041
rect 787 -1061 791 -1041
rect -356 -1144 -352 -1124
rect -348 -1144 -344 -1124
rect -304 -1144 -300 -1124
rect -296 -1144 -292 -1124
rect -460 -1191 -456 -1171
rect -452 -1191 -448 -1171
rect -408 -1191 -404 -1171
rect -400 -1191 -396 -1171
rect -356 -1191 -352 -1171
rect -348 -1191 -344 -1171
rect -304 -1191 -300 -1171
rect -296 -1191 -292 -1171
rect 593 -1345 597 -1305
rect 601 -1345 605 -1305
rect 593 -1410 597 -1370
rect 601 -1410 605 -1370
rect 636 -1379 640 -1359
rect 644 -1379 648 -1359
rect -268 -1448 -264 -1428
rect -260 -1448 -256 -1428
rect -236 -1448 -232 -1428
rect -228 -1448 -224 -1428
rect -365 -1472 -361 -1452
rect -357 -1472 -353 -1452
rect -313 -1472 -309 -1452
rect -305 -1472 -301 -1452
rect 80 -1487 100 -1483
rect 80 -1495 100 -1491
rect -469 -1519 -465 -1499
rect -461 -1519 -457 -1499
rect -417 -1519 -413 -1499
rect -409 -1519 -405 -1499
rect -365 -1519 -361 -1499
rect -357 -1519 -353 -1499
rect -313 -1519 -309 -1499
rect -305 -1519 -301 -1499
rect 178 -1502 182 -1482
rect 186 -1502 190 -1482
rect 80 -1538 100 -1534
rect 178 -1535 182 -1515
rect 186 -1535 190 -1515
rect 214 -1537 218 -1517
rect 222 -1537 226 -1517
rect 80 -1546 100 -1542
rect 594 -1628 598 -1588
rect 602 -1628 606 -1588
rect 830 -1575 834 -1535
rect 838 -1575 842 -1535
rect 1139 -1533 1143 -1513
rect 1147 -1533 1151 -1513
rect 1172 -1533 1176 -1513
rect 1180 -1533 1184 -1513
rect 1203 -1523 1207 -1503
rect 1211 -1523 1215 -1503
rect 830 -1640 834 -1600
rect 838 -1640 842 -1600
rect 873 -1609 877 -1589
rect 881 -1609 885 -1589
rect 150 -1717 154 -1677
rect 158 -1717 162 -1677
rect 594 -1693 598 -1653
rect 602 -1693 606 -1653
rect 637 -1662 641 -1642
rect 645 -1662 649 -1642
rect 150 -1782 154 -1742
rect 158 -1782 162 -1742
rect 193 -1751 197 -1731
rect 201 -1751 205 -1731
rect -284 -1826 -280 -1806
rect -276 -1826 -272 -1806
rect -252 -1826 -248 -1806
rect -244 -1826 -240 -1806
rect 839 -1786 843 -1746
rect 847 -1786 851 -1746
rect -381 -1850 -377 -1830
rect -373 -1850 -369 -1830
rect -329 -1850 -325 -1830
rect -321 -1850 -317 -1830
rect -485 -1897 -481 -1877
rect -477 -1897 -473 -1877
rect -433 -1897 -429 -1877
rect -425 -1897 -421 -1877
rect -381 -1897 -377 -1877
rect -373 -1897 -369 -1877
rect -329 -1897 -325 -1877
rect -321 -1897 -317 -1877
rect 590 -1899 594 -1859
rect 598 -1899 602 -1859
rect 839 -1851 843 -1811
rect 847 -1851 851 -1811
rect 882 -1820 886 -1800
rect 890 -1820 894 -1800
rect 1299 -1697 1303 -1677
rect 1307 -1697 1311 -1677
rect 1332 -1697 1336 -1677
rect 1340 -1697 1344 -1677
rect 1363 -1687 1367 -1667
rect 1371 -1687 1375 -1667
rect 1458 -1796 1478 -1792
rect 1150 -1833 1154 -1813
rect 1158 -1833 1162 -1813
rect 1183 -1833 1187 -1813
rect 1191 -1833 1195 -1813
rect 1214 -1823 1218 -1803
rect 1222 -1823 1226 -1803
rect 1458 -1804 1478 -1800
rect 1556 -1811 1560 -1791
rect 1564 -1811 1568 -1791
rect 1458 -1847 1478 -1843
rect 1556 -1844 1560 -1824
rect 1564 -1844 1568 -1824
rect 1592 -1846 1596 -1826
rect 1600 -1846 1604 -1826
rect 1458 -1855 1478 -1851
rect 2112 -1835 2116 -1815
rect 2120 -1835 2124 -1815
rect 2144 -1835 2148 -1815
rect 2152 -1835 2156 -1815
rect 2015 -1859 2019 -1839
rect 2023 -1859 2027 -1839
rect 2067 -1859 2071 -1839
rect 2075 -1859 2079 -1839
rect 1911 -1906 1915 -1886
rect 1919 -1906 1923 -1886
rect 1963 -1906 1967 -1886
rect 1971 -1906 1975 -1886
rect 2015 -1906 2019 -1886
rect 2023 -1906 2027 -1886
rect 2067 -1906 2071 -1886
rect 2075 -1906 2079 -1886
rect 590 -1964 594 -1924
rect 598 -1964 602 -1924
rect 633 -1933 637 -1913
rect 641 -1933 645 -1913
rect 578 -2148 582 -2108
rect 586 -2148 590 -2108
rect -268 -2196 -264 -2176
rect -260 -2196 -256 -2176
rect -236 -2196 -232 -2176
rect -228 -2196 -224 -2176
rect -365 -2220 -361 -2200
rect -357 -2220 -353 -2200
rect -313 -2220 -309 -2200
rect -305 -2220 -301 -2200
rect 578 -2213 582 -2173
rect 586 -2213 590 -2173
rect 621 -2182 625 -2162
rect 629 -2182 633 -2162
rect -469 -2267 -465 -2247
rect -461 -2267 -457 -2247
rect -417 -2267 -413 -2247
rect -409 -2267 -405 -2247
rect -365 -2267 -361 -2247
rect -357 -2267 -353 -2247
rect -313 -2267 -309 -2247
rect -305 -2267 -301 -2247
rect 77 -2362 97 -2358
rect 77 -2370 97 -2366
rect 175 -2377 179 -2357
rect 183 -2377 187 -2357
rect 77 -2413 97 -2409
rect 175 -2410 179 -2390
rect 183 -2410 187 -2390
rect 211 -2412 215 -2392
rect 219 -2412 223 -2392
rect 77 -2421 97 -2417
rect 717 -2458 721 -2418
rect 725 -2458 729 -2418
rect 717 -2523 721 -2483
rect 725 -2523 729 -2483
rect 760 -2492 764 -2472
rect 768 -2492 772 -2472
rect 1052 -2510 1056 -2470
rect 1060 -2510 1064 -2470
rect 147 -2592 151 -2552
rect 155 -2592 159 -2552
rect -259 -2625 -255 -2605
rect -251 -2625 -247 -2605
rect -227 -2625 -223 -2605
rect -219 -2625 -215 -2605
rect 1052 -2575 1056 -2535
rect 1060 -2575 1064 -2535
rect 1095 -2544 1099 -2524
rect 1103 -2544 1107 -2524
rect 1348 -2562 1352 -2542
rect 1356 -2562 1360 -2542
rect 1381 -2562 1385 -2542
rect 1389 -2562 1393 -2542
rect 1412 -2552 1416 -2532
rect 1420 -2552 1424 -2532
rect 2642 -2516 2646 -2496
rect 2650 -2516 2654 -2496
rect 2674 -2516 2678 -2496
rect 2682 -2516 2686 -2496
rect 2545 -2540 2549 -2520
rect 2553 -2540 2557 -2520
rect 2597 -2540 2601 -2520
rect 2605 -2540 2609 -2520
rect 2083 -2586 2087 -2566
rect 2091 -2586 2095 -2566
rect 2116 -2586 2120 -2566
rect 2124 -2586 2128 -2566
rect 2147 -2576 2151 -2556
rect 2155 -2576 2159 -2556
rect 2441 -2587 2445 -2567
rect 2449 -2587 2453 -2567
rect 2493 -2587 2497 -2567
rect 2501 -2587 2505 -2567
rect 2545 -2587 2549 -2567
rect 2553 -2587 2557 -2567
rect 2597 -2587 2601 -2567
rect 2605 -2587 2609 -2567
rect -356 -2649 -352 -2629
rect -348 -2649 -344 -2629
rect -304 -2649 -300 -2629
rect -296 -2649 -292 -2629
rect 147 -2657 151 -2617
rect 155 -2657 159 -2617
rect 190 -2626 194 -2606
rect 198 -2626 202 -2606
rect -460 -2696 -456 -2676
rect -452 -2696 -448 -2676
rect -408 -2696 -404 -2676
rect -400 -2696 -396 -2676
rect -356 -2696 -352 -2676
rect -348 -2696 -344 -2676
rect -304 -2696 -300 -2676
rect -296 -2696 -292 -2676
rect 718 -2741 722 -2701
rect 726 -2741 730 -2701
rect 718 -2806 722 -2766
rect 726 -2806 730 -2766
rect 761 -2775 765 -2755
rect 769 -2775 773 -2755
rect 1053 -2793 1057 -2753
rect 1061 -2793 1065 -2753
rect 1053 -2858 1057 -2818
rect 1061 -2858 1065 -2818
rect 1096 -2827 1100 -2807
rect 1104 -2827 1108 -2807
rect 1355 -2951 1359 -2931
rect 1363 -2951 1367 -2931
rect 1388 -2951 1392 -2931
rect 1396 -2951 1400 -2931
rect 1419 -2941 1423 -2921
rect 1427 -2941 1431 -2921
rect 714 -3012 718 -2972
rect 722 -3012 726 -2972
rect 714 -3077 718 -3037
rect 722 -3077 726 -3037
rect 757 -3046 761 -3026
rect 765 -3046 769 -3026
rect 1647 -3107 1651 -3087
rect 1655 -3107 1659 -3087
rect 1680 -3107 1684 -3087
rect 1688 -3107 1692 -3087
rect 1711 -3097 1715 -3077
rect 1719 -3097 1723 -3077
rect 1383 -3195 1387 -3155
rect 1391 -3195 1395 -3155
rect 702 -3261 706 -3221
rect 710 -3261 714 -3221
rect 702 -3326 706 -3286
rect 710 -3326 714 -3286
rect 745 -3295 749 -3275
rect 753 -3295 757 -3275
rect 1383 -3260 1387 -3220
rect 1391 -3260 1395 -3220
rect 1426 -3229 1430 -3209
rect 1434 -3229 1438 -3209
rect 1043 -3327 1047 -3287
rect 1051 -3327 1055 -3287
rect 1043 -3392 1047 -3352
rect 1051 -3392 1055 -3352
rect 1086 -3361 1090 -3341
rect 1094 -3361 1098 -3341
rect 719 -3528 723 -3488
rect 727 -3528 731 -3488
rect 719 -3593 723 -3553
rect 727 -3593 731 -3553
rect 762 -3562 766 -3542
rect 770 -3562 774 -3542
rect 707 -3777 711 -3737
rect 715 -3777 719 -3737
rect 707 -3842 711 -3802
rect 715 -3842 719 -3802
rect 750 -3811 754 -3791
rect 758 -3811 762 -3791
<< pdcontact >>
rect 1171 165 1175 205
rect 1179 165 1183 205
rect 1223 165 1227 205
rect 1231 165 1235 205
rect 1275 165 1279 205
rect 1283 165 1287 205
rect 1327 165 1331 205
rect 1335 165 1339 205
rect 1372 173 1376 213
rect 1380 173 1384 213
rect 1404 173 1408 213
rect 1412 173 1416 213
rect 1171 103 1175 143
rect 1179 103 1183 143
rect 1223 103 1227 143
rect 1231 103 1235 143
rect -460 39 -456 79
rect -452 39 -448 79
rect -408 39 -404 79
rect -400 39 -396 79
rect -356 39 -352 79
rect -348 39 -344 79
rect -304 39 -300 79
rect -296 39 -292 79
rect -259 47 -255 87
rect -251 47 -247 87
rect -227 47 -223 87
rect -219 47 -215 87
rect -460 -23 -456 17
rect -452 -23 -448 17
rect -408 -23 -404 17
rect -400 -23 -396 17
rect 530 0 570 4
rect 530 -8 570 -4
rect 626 -12 630 28
rect 634 -12 638 28
rect 530 -51 570 -47
rect 530 -59 570 -55
rect 158 -191 198 -187
rect 158 -199 198 -195
rect 254 -203 258 -163
rect 262 -203 266 -163
rect 158 -242 198 -238
rect 475 -219 479 -179
rect 483 -219 487 -179
rect 502 -219 506 -179
rect 510 -219 514 -179
rect 158 -250 198 -246
rect 720 -226 724 -146
rect 728 -226 732 -146
rect -427 -356 -423 -316
rect -419 -356 -415 -316
rect -375 -356 -371 -316
rect -367 -356 -363 -316
rect -323 -356 -319 -316
rect -315 -356 -311 -316
rect -271 -356 -267 -316
rect -263 -356 -259 -316
rect -226 -348 -222 -308
rect -218 -348 -214 -308
rect -194 -348 -190 -308
rect -186 -348 -182 -308
rect 171 -347 175 -307
rect 179 -347 183 -307
rect 198 -347 202 -307
rect 206 -347 210 -307
rect 537 -289 541 -249
rect 545 -289 549 -249
rect -427 -418 -423 -378
rect -419 -418 -415 -378
rect -375 -418 -371 -378
rect -367 -418 -363 -378
rect 720 -326 724 -246
rect 728 -326 732 -246
rect 769 -323 773 -283
rect 777 -323 781 -283
rect 1449 -298 1453 -258
rect 1457 -298 1461 -258
rect 1501 -298 1505 -258
rect 1509 -298 1513 -258
rect 1553 -298 1557 -258
rect 1561 -298 1565 -258
rect 1605 -298 1609 -258
rect 1613 -298 1617 -258
rect 1650 -290 1654 -250
rect 1658 -290 1662 -250
rect 1682 -290 1686 -250
rect 1690 -290 1694 -250
rect 233 -417 237 -377
rect 241 -417 245 -377
rect 1026 -387 1066 -383
rect 1026 -395 1066 -391
rect 1122 -399 1126 -359
rect 1130 -399 1134 -359
rect 1449 -360 1453 -320
rect 1457 -360 1461 -320
rect 1501 -360 1505 -320
rect 1509 -360 1513 -320
rect 1026 -438 1066 -434
rect 1026 -446 1066 -442
rect -536 -735 -532 -695
rect -528 -735 -524 -695
rect -484 -735 -480 -695
rect -476 -735 -472 -695
rect -432 -735 -428 -695
rect -424 -735 -420 -695
rect -380 -735 -376 -695
rect -372 -735 -368 -695
rect -335 -727 -331 -687
rect -327 -727 -323 -687
rect -303 -727 -299 -687
rect -295 -727 -291 -687
rect 576 -708 580 -668
rect 584 -708 588 -668
rect 603 -708 607 -668
rect 611 -708 615 -668
rect 975 -715 979 -635
rect 983 -715 987 -635
rect 1201 -707 1205 -627
rect 1209 -707 1213 -627
rect -536 -797 -532 -757
rect -528 -797 -524 -757
rect -484 -797 -480 -757
rect -476 -797 -472 -757
rect 638 -778 642 -738
rect 646 -778 650 -738
rect 109 -827 149 -823
rect 109 -835 149 -831
rect 205 -839 209 -799
rect 213 -839 217 -799
rect 109 -878 149 -874
rect 975 -815 979 -735
rect 983 -815 987 -735
rect 1024 -812 1028 -772
rect 1032 -812 1036 -772
rect 1201 -807 1205 -727
rect 1209 -807 1213 -727
rect 1250 -804 1254 -764
rect 1258 -804 1262 -764
rect 1380 -832 1420 -828
rect 1380 -840 1420 -836
rect 1476 -844 1480 -804
rect 1484 -844 1488 -804
rect 109 -886 149 -882
rect 1380 -883 1420 -879
rect 1760 -853 1764 -813
rect 1768 -853 1772 -813
rect 1812 -853 1816 -813
rect 1820 -853 1824 -813
rect 1864 -853 1868 -813
rect 1872 -853 1876 -813
rect 1916 -853 1920 -813
rect 1924 -853 1928 -813
rect 1961 -845 1965 -805
rect 1969 -845 1973 -805
rect 1993 -845 1997 -805
rect 2001 -845 2005 -805
rect 1380 -891 1420 -887
rect 122 -983 126 -943
rect 130 -983 134 -943
rect 149 -983 153 -943
rect 157 -983 161 -943
rect 499 -953 503 -913
rect 507 -953 511 -913
rect 526 -953 530 -913
rect 534 -953 538 -913
rect 717 -953 721 -913
rect 725 -953 729 -913
rect 744 -953 748 -913
rect 752 -953 756 -913
rect 1760 -915 1764 -875
rect 1768 -915 1772 -875
rect 1812 -915 1816 -875
rect 1820 -915 1824 -875
rect -460 -1088 -456 -1048
rect -452 -1088 -448 -1048
rect -408 -1088 -404 -1048
rect -400 -1088 -396 -1048
rect -356 -1088 -352 -1048
rect -348 -1088 -344 -1048
rect -304 -1088 -300 -1048
rect -296 -1088 -292 -1048
rect -259 -1080 -255 -1040
rect -251 -1080 -247 -1040
rect -227 -1080 -223 -1040
rect -219 -1080 -215 -1040
rect 184 -1053 188 -1013
rect 192 -1053 196 -1013
rect 561 -1023 565 -983
rect 569 -1023 573 -983
rect -460 -1150 -456 -1110
rect -452 -1150 -448 -1110
rect -408 -1150 -404 -1110
rect -400 -1150 -396 -1110
rect 779 -1023 783 -983
rect 787 -1023 791 -983
rect 574 -1271 578 -1231
rect 582 -1271 586 -1231
rect 601 -1271 605 -1231
rect 609 -1271 613 -1231
rect 636 -1341 640 -1301
rect 644 -1341 648 -1301
rect -469 -1416 -465 -1376
rect -461 -1416 -457 -1376
rect -417 -1416 -413 -1376
rect -409 -1416 -405 -1376
rect -365 -1416 -361 -1376
rect -357 -1416 -353 -1376
rect -313 -1416 -309 -1376
rect -305 -1416 -301 -1376
rect -268 -1408 -264 -1368
rect -260 -1408 -256 -1368
rect -236 -1408 -232 -1368
rect -228 -1408 -224 -1368
rect 1154 -1388 1158 -1308
rect 1162 -1388 1166 -1308
rect -469 -1478 -465 -1438
rect -461 -1478 -457 -1438
rect -417 -1478 -413 -1438
rect -409 -1478 -405 -1438
rect 118 -1487 158 -1483
rect 118 -1495 158 -1491
rect 214 -1499 218 -1459
rect 222 -1499 226 -1459
rect 118 -1538 158 -1534
rect 811 -1501 815 -1461
rect 819 -1501 823 -1461
rect 838 -1501 842 -1461
rect 846 -1501 850 -1461
rect 1154 -1488 1158 -1408
rect 1162 -1488 1166 -1408
rect 118 -1546 158 -1542
rect 575 -1554 579 -1514
rect 583 -1554 587 -1514
rect 602 -1554 606 -1514
rect 610 -1554 614 -1514
rect 1203 -1485 1207 -1445
rect 1211 -1485 1215 -1445
rect 131 -1643 135 -1603
rect 139 -1643 143 -1603
rect 158 -1643 162 -1603
rect 166 -1643 170 -1603
rect 637 -1624 641 -1584
rect 645 -1624 649 -1584
rect 873 -1571 877 -1531
rect 881 -1571 885 -1531
rect 1314 -1552 1318 -1472
rect 1322 -1552 1326 -1472
rect 193 -1713 197 -1673
rect 201 -1713 205 -1673
rect 820 -1712 824 -1672
rect 828 -1712 832 -1672
rect 847 -1712 851 -1672
rect 855 -1712 859 -1672
rect 1165 -1688 1169 -1608
rect 1173 -1688 1177 -1608
rect 1314 -1652 1318 -1572
rect 1322 -1652 1326 -1572
rect 1363 -1649 1367 -1609
rect 1371 -1649 1375 -1609
rect -485 -1794 -481 -1754
rect -477 -1794 -473 -1754
rect -433 -1794 -429 -1754
rect -425 -1794 -421 -1754
rect -381 -1794 -377 -1754
rect -373 -1794 -369 -1754
rect -329 -1794 -325 -1754
rect -321 -1794 -317 -1754
rect -284 -1786 -280 -1746
rect -276 -1786 -272 -1746
rect -252 -1786 -248 -1746
rect -244 -1786 -240 -1746
rect -485 -1856 -481 -1816
rect -477 -1856 -473 -1816
rect -433 -1856 -429 -1816
rect -425 -1856 -421 -1816
rect 571 -1825 575 -1785
rect 579 -1825 583 -1785
rect 598 -1825 602 -1785
rect 606 -1825 610 -1785
rect 882 -1782 886 -1742
rect 890 -1782 894 -1742
rect 1165 -1788 1169 -1708
rect 1173 -1788 1177 -1708
rect 1214 -1785 1218 -1745
rect 1222 -1785 1226 -1745
rect 1496 -1796 1536 -1792
rect 1496 -1804 1536 -1800
rect 1592 -1808 1596 -1768
rect 1600 -1808 1604 -1768
rect 1911 -1803 1915 -1763
rect 1919 -1803 1923 -1763
rect 1963 -1803 1967 -1763
rect 1971 -1803 1975 -1763
rect 2015 -1803 2019 -1763
rect 2023 -1803 2027 -1763
rect 2067 -1803 2071 -1763
rect 2075 -1803 2079 -1763
rect 2112 -1795 2116 -1755
rect 2120 -1795 2124 -1755
rect 2144 -1795 2148 -1755
rect 2152 -1795 2156 -1755
rect 1496 -1847 1536 -1843
rect 1496 -1855 1536 -1851
rect 633 -1895 637 -1855
rect 641 -1895 645 -1855
rect 1911 -1865 1915 -1825
rect 1919 -1865 1923 -1825
rect 1963 -1865 1967 -1825
rect 1971 -1865 1975 -1825
rect 559 -2074 563 -2034
rect 567 -2074 571 -2034
rect 586 -2074 590 -2034
rect 594 -2074 598 -2034
rect -469 -2164 -465 -2124
rect -461 -2164 -457 -2124
rect -417 -2164 -413 -2124
rect -409 -2164 -405 -2124
rect -365 -2164 -361 -2124
rect -357 -2164 -353 -2124
rect -313 -2164 -309 -2124
rect -305 -2164 -301 -2124
rect -268 -2156 -264 -2116
rect -260 -2156 -256 -2116
rect -236 -2156 -232 -2116
rect -228 -2156 -224 -2116
rect 621 -2144 625 -2104
rect 629 -2144 633 -2104
rect -469 -2226 -465 -2186
rect -461 -2226 -457 -2186
rect -417 -2226 -413 -2186
rect -409 -2226 -405 -2186
rect 115 -2362 155 -2358
rect 115 -2370 155 -2366
rect 211 -2374 215 -2334
rect 219 -2374 223 -2334
rect 115 -2413 155 -2409
rect 698 -2384 702 -2344
rect 706 -2384 710 -2344
rect 725 -2384 729 -2344
rect 733 -2384 737 -2344
rect 115 -2421 155 -2417
rect 760 -2454 764 -2414
rect 768 -2454 772 -2414
rect 1033 -2436 1037 -2396
rect 1041 -2436 1045 -2396
rect 1060 -2436 1064 -2396
rect 1068 -2436 1072 -2396
rect 1363 -2417 1367 -2337
rect 1371 -2417 1375 -2337
rect 128 -2518 132 -2478
rect 136 -2518 140 -2478
rect 155 -2518 159 -2478
rect 163 -2518 167 -2478
rect -460 -2593 -456 -2553
rect -452 -2593 -448 -2553
rect -408 -2593 -404 -2553
rect -400 -2593 -396 -2553
rect -356 -2593 -352 -2553
rect -348 -2593 -344 -2553
rect -304 -2593 -300 -2553
rect -296 -2593 -292 -2553
rect -259 -2585 -255 -2545
rect -251 -2585 -247 -2545
rect -227 -2585 -223 -2545
rect -219 -2585 -215 -2545
rect 1095 -2506 1099 -2466
rect 1103 -2506 1107 -2466
rect 1363 -2517 1367 -2437
rect 1371 -2517 1375 -2437
rect -460 -2655 -456 -2615
rect -452 -2655 -448 -2615
rect -408 -2655 -404 -2615
rect -400 -2655 -396 -2615
rect 190 -2588 194 -2548
rect 198 -2588 202 -2548
rect 2098 -2441 2102 -2361
rect 2106 -2441 2110 -2361
rect 1412 -2514 1416 -2474
rect 1420 -2514 1424 -2474
rect 2098 -2541 2102 -2461
rect 2106 -2541 2110 -2461
rect 2441 -2484 2445 -2444
rect 2449 -2484 2453 -2444
rect 2493 -2484 2497 -2444
rect 2501 -2484 2505 -2444
rect 2545 -2484 2549 -2444
rect 2553 -2484 2557 -2444
rect 2597 -2484 2601 -2444
rect 2605 -2484 2609 -2444
rect 2642 -2476 2646 -2436
rect 2650 -2476 2654 -2436
rect 2674 -2476 2678 -2436
rect 2682 -2476 2686 -2436
rect 2147 -2538 2151 -2498
rect 2155 -2538 2159 -2498
rect 2441 -2546 2445 -2506
rect 2449 -2546 2453 -2506
rect 2493 -2546 2497 -2506
rect 2501 -2546 2505 -2506
rect 699 -2667 703 -2627
rect 707 -2667 711 -2627
rect 726 -2667 730 -2627
rect 734 -2667 738 -2627
rect 761 -2737 765 -2697
rect 769 -2737 773 -2697
rect 1034 -2719 1038 -2679
rect 1042 -2719 1046 -2679
rect 1061 -2719 1065 -2679
rect 1069 -2719 1073 -2679
rect 1096 -2789 1100 -2749
rect 1104 -2789 1108 -2749
rect 1370 -2806 1374 -2726
rect 1378 -2806 1382 -2726
rect 695 -2938 699 -2898
rect 703 -2938 707 -2898
rect 722 -2938 726 -2898
rect 730 -2938 734 -2898
rect 1370 -2906 1374 -2826
rect 1378 -2906 1382 -2826
rect 1419 -2903 1423 -2863
rect 1427 -2903 1431 -2863
rect 1662 -2962 1666 -2882
rect 1670 -2962 1674 -2882
rect 757 -3008 761 -2968
rect 765 -3008 769 -2968
rect 1662 -3062 1666 -2982
rect 1670 -3062 1674 -2982
rect 1364 -3121 1368 -3081
rect 1372 -3121 1376 -3081
rect 1391 -3121 1395 -3081
rect 1399 -3121 1403 -3081
rect 1711 -3059 1715 -3019
rect 1719 -3059 1723 -3019
rect 683 -3187 687 -3147
rect 691 -3187 695 -3147
rect 710 -3187 714 -3147
rect 718 -3187 722 -3147
rect 1426 -3191 1430 -3151
rect 1434 -3191 1438 -3151
rect 745 -3257 749 -3217
rect 753 -3257 757 -3217
rect 1024 -3253 1028 -3213
rect 1032 -3253 1036 -3213
rect 1051 -3253 1055 -3213
rect 1059 -3253 1063 -3213
rect 1086 -3323 1090 -3283
rect 1094 -3323 1098 -3283
rect 700 -3454 704 -3414
rect 708 -3454 712 -3414
rect 727 -3454 731 -3414
rect 735 -3454 739 -3414
rect 762 -3524 766 -3484
rect 770 -3524 774 -3484
rect 688 -3703 692 -3663
rect 696 -3703 700 -3663
rect 715 -3703 719 -3663
rect 723 -3703 727 -3663
rect 750 -3773 754 -3733
rect 758 -3773 762 -3733
<< psubstratepcontact >>
rect 1364 120 1368 124
rect 1388 120 1392 124
rect 1396 120 1400 124
rect 1420 120 1424 124
rect 1188 49 1192 53
rect 1240 49 1244 53
rect 1292 49 1296 53
rect 1344 49 1348 53
rect 481 7 485 11
rect -267 -6 -263 -2
rect -243 -6 -239 -2
rect -235 -6 -231 -2
rect -211 -6 -207 -2
rect 481 -14 485 -10
rect 481 -44 485 -40
rect 481 -65 485 -61
rect 619 -61 623 -57
rect 640 -61 644 -57
rect -443 -77 -439 -73
rect -391 -77 -387 -73
rect -339 -77 -335 -73
rect -287 -77 -283 -73
rect 109 -184 113 -180
rect 109 -205 113 -201
rect 109 -235 113 -231
rect 109 -256 113 -252
rect 247 -252 251 -248
rect 268 -252 272 -248
rect 530 -338 534 -334
rect 551 -338 555 -334
rect -234 -401 -230 -397
rect -210 -401 -206 -397
rect -202 -401 -198 -397
rect -178 -401 -174 -397
rect 487 -369 491 -365
rect 508 -369 512 -365
rect 762 -372 766 -368
rect 783 -372 787 -368
rect 698 -382 702 -378
rect 719 -382 723 -378
rect 731 -382 735 -378
rect 752 -382 756 -378
rect 977 -380 981 -376
rect 977 -401 981 -397
rect 1642 -343 1646 -339
rect 1666 -343 1670 -339
rect 1674 -343 1678 -339
rect 1698 -343 1702 -339
rect 977 -431 981 -427
rect -410 -472 -406 -468
rect -358 -472 -354 -468
rect -306 -472 -302 -468
rect -254 -472 -250 -468
rect 1466 -414 1470 -410
rect 1518 -414 1522 -410
rect 1570 -414 1574 -410
rect 1622 -414 1626 -410
rect 977 -452 981 -448
rect 1115 -448 1119 -444
rect 1136 -448 1140 -444
rect 226 -466 230 -462
rect 247 -466 251 -462
rect 183 -497 187 -493
rect 204 -497 208 -493
rect -343 -780 -339 -776
rect -319 -780 -315 -776
rect -311 -780 -307 -776
rect -287 -780 -283 -776
rect 60 -820 64 -816
rect 60 -841 64 -837
rect -519 -851 -515 -847
rect -467 -851 -463 -847
rect -415 -851 -411 -847
rect -363 -851 -359 -847
rect 60 -871 64 -867
rect 631 -827 635 -823
rect 652 -827 656 -823
rect 588 -858 592 -854
rect 609 -858 613 -854
rect 1331 -825 1335 -821
rect 1331 -846 1335 -842
rect 1243 -853 1247 -849
rect 1264 -853 1268 -849
rect 1017 -861 1021 -857
rect 1038 -861 1042 -857
rect 1179 -863 1183 -859
rect 1200 -863 1204 -859
rect 1212 -863 1216 -859
rect 1233 -863 1237 -859
rect 953 -871 957 -867
rect 974 -871 978 -867
rect 986 -871 990 -867
rect 1007 -871 1011 -867
rect 1331 -876 1335 -872
rect 60 -892 64 -888
rect 198 -888 202 -884
rect 219 -888 223 -884
rect 1331 -897 1335 -893
rect 1469 -893 1473 -889
rect 1490 -893 1494 -889
rect 1953 -898 1957 -894
rect 1977 -898 1981 -894
rect 1985 -898 1989 -894
rect 2009 -898 2013 -894
rect 1777 -969 1781 -965
rect 1829 -969 1833 -965
rect 1881 -969 1885 -965
rect 1933 -969 1937 -965
rect 554 -1072 558 -1068
rect 575 -1072 579 -1068
rect 772 -1072 776 -1068
rect 793 -1072 797 -1068
rect 177 -1102 181 -1098
rect 198 -1102 202 -1098
rect 511 -1103 515 -1099
rect 532 -1103 536 -1099
rect 729 -1103 733 -1099
rect 750 -1103 754 -1099
rect -267 -1133 -263 -1129
rect -243 -1133 -239 -1129
rect -235 -1133 -231 -1129
rect -211 -1133 -207 -1129
rect 134 -1133 138 -1129
rect 155 -1133 159 -1129
rect -443 -1204 -439 -1200
rect -391 -1204 -387 -1200
rect -339 -1204 -335 -1200
rect -287 -1204 -283 -1200
rect 629 -1390 633 -1386
rect 650 -1390 654 -1386
rect 586 -1421 590 -1417
rect 607 -1421 611 -1417
rect -276 -1461 -272 -1457
rect -252 -1461 -248 -1457
rect -244 -1461 -240 -1457
rect -220 -1461 -216 -1457
rect 69 -1480 73 -1476
rect 69 -1501 73 -1497
rect -452 -1532 -448 -1528
rect -400 -1532 -396 -1528
rect -348 -1532 -344 -1528
rect -296 -1532 -292 -1528
rect 69 -1531 73 -1527
rect 69 -1552 73 -1548
rect 207 -1548 211 -1544
rect 228 -1548 232 -1544
rect 1196 -1534 1200 -1530
rect 1217 -1534 1221 -1530
rect 1132 -1544 1136 -1540
rect 1153 -1544 1157 -1540
rect 1165 -1544 1169 -1540
rect 1186 -1544 1190 -1540
rect 866 -1620 870 -1616
rect 887 -1620 891 -1616
rect 823 -1651 827 -1647
rect 844 -1651 848 -1647
rect 630 -1673 634 -1669
rect 651 -1673 655 -1669
rect 587 -1704 591 -1700
rect 608 -1704 612 -1700
rect 186 -1762 190 -1758
rect 207 -1762 211 -1758
rect 143 -1793 147 -1789
rect 164 -1793 168 -1789
rect -292 -1839 -288 -1835
rect -268 -1839 -264 -1835
rect -260 -1839 -256 -1835
rect -236 -1839 -232 -1835
rect -468 -1910 -464 -1906
rect -416 -1910 -412 -1906
rect -364 -1910 -360 -1906
rect -312 -1910 -308 -1906
rect 1356 -1698 1360 -1694
rect 1377 -1698 1381 -1694
rect 1292 -1708 1296 -1704
rect 1313 -1708 1317 -1704
rect 1325 -1708 1329 -1704
rect 1346 -1708 1350 -1704
rect 1447 -1789 1451 -1785
rect 875 -1831 879 -1827
rect 896 -1831 900 -1827
rect 1447 -1810 1451 -1806
rect 1207 -1834 1211 -1830
rect 1228 -1834 1232 -1830
rect 1447 -1840 1451 -1836
rect 1143 -1844 1147 -1840
rect 1164 -1844 1168 -1840
rect 1176 -1844 1180 -1840
rect 1197 -1844 1201 -1840
rect 832 -1862 836 -1858
rect 853 -1862 857 -1858
rect 1447 -1861 1451 -1857
rect 1585 -1857 1589 -1853
rect 1606 -1857 1610 -1853
rect 2104 -1848 2108 -1844
rect 2128 -1848 2132 -1844
rect 2136 -1848 2140 -1844
rect 2160 -1848 2164 -1844
rect 1928 -1919 1932 -1915
rect 1980 -1919 1984 -1915
rect 2032 -1919 2036 -1915
rect 2084 -1919 2088 -1915
rect 626 -1944 630 -1940
rect 647 -1944 651 -1940
rect 583 -1975 587 -1971
rect 604 -1975 608 -1971
rect -276 -2209 -272 -2205
rect -252 -2209 -248 -2205
rect -244 -2209 -240 -2205
rect -220 -2209 -216 -2205
rect 614 -2193 618 -2189
rect 635 -2193 639 -2189
rect 571 -2224 575 -2220
rect 592 -2224 596 -2220
rect -452 -2280 -448 -2276
rect -400 -2280 -396 -2276
rect -348 -2280 -344 -2276
rect -296 -2280 -292 -2276
rect 66 -2355 70 -2351
rect 66 -2376 70 -2372
rect 66 -2406 70 -2402
rect 66 -2427 70 -2423
rect 204 -2423 208 -2419
rect 225 -2423 229 -2419
rect 753 -2503 757 -2499
rect 774 -2503 778 -2499
rect 710 -2534 714 -2530
rect 731 -2534 735 -2530
rect 1088 -2555 1092 -2551
rect 1109 -2555 1113 -2551
rect 1405 -2563 1409 -2559
rect 1426 -2563 1430 -2559
rect 2634 -2529 2638 -2525
rect 2658 -2529 2662 -2525
rect 2666 -2529 2670 -2525
rect 2690 -2529 2694 -2525
rect 1341 -2573 1345 -2569
rect 1362 -2573 1366 -2569
rect 1374 -2573 1378 -2569
rect 1395 -2573 1399 -2569
rect 1045 -2586 1049 -2582
rect 1066 -2586 1070 -2582
rect 2140 -2587 2144 -2583
rect 2161 -2587 2165 -2583
rect 2076 -2597 2080 -2593
rect 2097 -2597 2101 -2593
rect 2109 -2597 2113 -2593
rect 2130 -2597 2134 -2593
rect 2458 -2600 2462 -2596
rect 2510 -2600 2514 -2596
rect 2562 -2600 2566 -2596
rect 2614 -2600 2618 -2596
rect -267 -2638 -263 -2634
rect -243 -2638 -239 -2634
rect -235 -2638 -231 -2634
rect -211 -2638 -207 -2634
rect 183 -2637 187 -2633
rect 204 -2637 208 -2633
rect 140 -2668 144 -2664
rect 161 -2668 165 -2664
rect -443 -2709 -439 -2705
rect -391 -2709 -387 -2705
rect -339 -2709 -335 -2705
rect -287 -2709 -283 -2705
rect 754 -2786 758 -2782
rect 775 -2786 779 -2782
rect 711 -2817 715 -2813
rect 732 -2817 736 -2813
rect 1089 -2838 1093 -2834
rect 1110 -2838 1114 -2834
rect 1046 -2869 1050 -2865
rect 1067 -2869 1071 -2865
rect 1412 -2952 1416 -2948
rect 1433 -2952 1437 -2948
rect 1348 -2962 1352 -2958
rect 1369 -2962 1373 -2958
rect 1381 -2962 1385 -2958
rect 1402 -2962 1406 -2958
rect 750 -3057 754 -3053
rect 771 -3057 775 -3053
rect 707 -3088 711 -3084
rect 728 -3088 732 -3084
rect 1704 -3108 1708 -3104
rect 1725 -3108 1729 -3104
rect 1640 -3118 1644 -3114
rect 1661 -3118 1665 -3114
rect 1673 -3118 1677 -3114
rect 1694 -3118 1698 -3114
rect 1419 -3240 1423 -3236
rect 1440 -3240 1444 -3236
rect 738 -3306 742 -3302
rect 759 -3306 763 -3302
rect 695 -3337 699 -3333
rect 716 -3337 720 -3333
rect 1376 -3271 1380 -3267
rect 1397 -3271 1401 -3267
rect 1079 -3372 1083 -3368
rect 1100 -3372 1104 -3368
rect 1036 -3403 1040 -3399
rect 1057 -3403 1061 -3399
rect 755 -3573 759 -3569
rect 776 -3573 780 -3569
rect 712 -3604 716 -3600
rect 733 -3604 737 -3600
rect 743 -3822 747 -3818
rect 764 -3822 768 -3818
rect 700 -3853 704 -3849
rect 721 -3853 725 -3849
<< nsubstratencontact >>
rect 1365 221 1369 225
rect 1387 221 1391 225
rect 1397 221 1401 225
rect 1419 221 1423 225
rect 1164 213 1168 217
rect 1186 213 1190 217
rect 1216 213 1220 217
rect 1238 213 1242 217
rect 1268 213 1272 217
rect 1290 213 1294 217
rect 1320 213 1324 217
rect 1342 213 1346 217
rect -266 95 -262 99
rect -244 95 -240 99
rect -234 95 -230 99
rect -212 95 -208 99
rect -467 87 -463 91
rect -445 87 -441 91
rect -415 87 -411 91
rect -393 87 -389 91
rect -363 87 -359 91
rect -341 87 -337 91
rect -311 87 -307 91
rect -289 87 -285 91
rect 621 35 625 39
rect 638 35 642 39
rect 577 5 581 9
rect 577 -12 581 -8
rect 577 -46 581 -42
rect 577 -63 581 -59
rect 715 -139 719 -135
rect 732 -139 736 -135
rect 249 -156 253 -152
rect 266 -156 270 -152
rect 205 -186 209 -182
rect 205 -203 209 -199
rect 470 -172 474 -168
rect 487 -172 491 -168
rect 497 -172 501 -168
rect 514 -172 518 -168
rect 205 -237 209 -233
rect 205 -254 209 -250
rect -233 -300 -229 -296
rect -211 -300 -207 -296
rect -201 -300 -197 -296
rect -179 -300 -175 -296
rect 166 -300 170 -296
rect 183 -300 187 -296
rect 193 -300 197 -296
rect 210 -300 214 -296
rect -434 -308 -430 -304
rect -412 -308 -408 -304
rect -382 -308 -378 -304
rect -360 -308 -356 -304
rect -330 -308 -326 -304
rect -308 -308 -304 -304
rect -278 -308 -274 -304
rect -256 -308 -252 -304
rect 532 -242 536 -238
rect 549 -242 553 -238
rect 1643 -242 1647 -238
rect 1665 -242 1669 -238
rect 1675 -242 1679 -238
rect 1697 -242 1701 -238
rect 1442 -250 1446 -246
rect 1464 -250 1468 -246
rect 1494 -250 1498 -246
rect 1516 -250 1520 -246
rect 1546 -250 1550 -246
rect 1568 -250 1572 -246
rect 1598 -250 1602 -246
rect 1620 -250 1624 -246
rect 764 -276 768 -272
rect 781 -276 785 -272
rect 228 -370 232 -366
rect 245 -370 249 -366
rect 1117 -352 1121 -348
rect 1134 -352 1138 -348
rect 1073 -382 1077 -378
rect 1073 -399 1077 -395
rect 1073 -433 1077 -429
rect 1073 -450 1077 -446
rect 1196 -620 1200 -616
rect 1213 -620 1217 -616
rect 970 -628 974 -624
rect 987 -628 991 -624
rect 571 -661 575 -657
rect 588 -661 592 -657
rect 598 -661 602 -657
rect 615 -661 619 -657
rect -342 -679 -338 -675
rect -320 -679 -316 -675
rect -310 -679 -306 -675
rect -288 -679 -284 -675
rect -543 -687 -539 -683
rect -521 -687 -517 -683
rect -491 -687 -487 -683
rect -469 -687 -465 -683
rect -439 -687 -435 -683
rect -417 -687 -413 -683
rect -387 -687 -383 -683
rect -365 -687 -361 -683
rect 200 -792 204 -788
rect 217 -792 221 -788
rect 633 -731 637 -727
rect 650 -731 654 -727
rect 156 -822 160 -818
rect 156 -839 160 -835
rect 156 -873 160 -869
rect 1019 -765 1023 -761
rect 1036 -765 1040 -761
rect 1245 -757 1249 -753
rect 1262 -757 1266 -753
rect 1471 -797 1475 -793
rect 1488 -797 1492 -793
rect 1954 -797 1958 -793
rect 1976 -797 1980 -793
rect 1986 -797 1990 -793
rect 2008 -797 2012 -793
rect 1427 -827 1431 -823
rect 1427 -844 1431 -840
rect 1753 -805 1757 -801
rect 1775 -805 1779 -801
rect 1805 -805 1809 -801
rect 1827 -805 1831 -801
rect 1857 -805 1861 -801
rect 1879 -805 1883 -801
rect 1909 -805 1913 -801
rect 1931 -805 1935 -801
rect 1427 -878 1431 -874
rect 156 -890 160 -886
rect 1427 -895 1431 -891
rect 494 -906 498 -902
rect 511 -906 515 -902
rect 521 -906 525 -902
rect 538 -906 542 -902
rect 712 -906 716 -902
rect 729 -906 733 -902
rect 739 -906 743 -902
rect 756 -906 760 -902
rect 117 -936 121 -932
rect 134 -936 138 -932
rect 144 -936 148 -932
rect 161 -936 165 -932
rect -266 -1032 -262 -1028
rect -244 -1032 -240 -1028
rect -234 -1032 -230 -1028
rect -212 -1032 -208 -1028
rect -467 -1040 -463 -1036
rect -445 -1040 -441 -1036
rect -415 -1040 -411 -1036
rect -393 -1040 -389 -1036
rect -363 -1040 -359 -1036
rect -341 -1040 -337 -1036
rect -311 -1040 -307 -1036
rect -289 -1040 -285 -1036
rect 179 -1006 183 -1002
rect 196 -1006 200 -1002
rect 556 -976 560 -972
rect 573 -976 577 -972
rect 774 -976 778 -972
rect 791 -976 795 -972
rect 569 -1224 573 -1220
rect 586 -1224 590 -1220
rect 596 -1224 600 -1220
rect 613 -1224 617 -1220
rect -275 -1360 -271 -1356
rect -253 -1360 -249 -1356
rect -243 -1360 -239 -1356
rect -221 -1360 -217 -1356
rect 631 -1294 635 -1290
rect 648 -1294 652 -1290
rect 1149 -1301 1153 -1297
rect 1166 -1301 1170 -1297
rect -476 -1368 -472 -1364
rect -454 -1368 -450 -1364
rect -424 -1368 -420 -1364
rect -402 -1368 -398 -1364
rect -372 -1368 -368 -1364
rect -350 -1368 -346 -1364
rect -320 -1368 -316 -1364
rect -298 -1368 -294 -1364
rect 209 -1452 213 -1448
rect 226 -1452 230 -1448
rect 806 -1454 810 -1450
rect 823 -1454 827 -1450
rect 833 -1454 837 -1450
rect 850 -1454 854 -1450
rect 165 -1482 169 -1478
rect 165 -1499 169 -1495
rect 165 -1533 169 -1529
rect 570 -1507 574 -1503
rect 587 -1507 591 -1503
rect 597 -1507 601 -1503
rect 614 -1507 618 -1503
rect 165 -1550 169 -1546
rect 1198 -1438 1202 -1434
rect 1215 -1438 1219 -1434
rect 1309 -1465 1313 -1461
rect 1326 -1465 1330 -1461
rect 126 -1596 130 -1592
rect 143 -1596 147 -1592
rect 153 -1596 157 -1592
rect 170 -1596 174 -1592
rect 632 -1577 636 -1573
rect 649 -1577 653 -1573
rect 868 -1524 872 -1520
rect 885 -1524 889 -1520
rect 1160 -1601 1164 -1597
rect 1177 -1601 1181 -1597
rect 188 -1666 192 -1662
rect 205 -1666 209 -1662
rect 815 -1665 819 -1661
rect 832 -1665 836 -1661
rect 842 -1665 846 -1661
rect 859 -1665 863 -1661
rect 1358 -1602 1362 -1598
rect 1375 -1602 1379 -1598
rect -291 -1738 -287 -1734
rect -269 -1738 -265 -1734
rect -259 -1738 -255 -1734
rect -237 -1738 -233 -1734
rect -492 -1746 -488 -1742
rect -470 -1746 -466 -1742
rect -440 -1746 -436 -1742
rect -418 -1746 -414 -1742
rect -388 -1746 -384 -1742
rect -366 -1746 -362 -1742
rect -336 -1746 -332 -1742
rect -314 -1746 -310 -1742
rect 566 -1778 570 -1774
rect 583 -1778 587 -1774
rect 593 -1778 597 -1774
rect 610 -1778 614 -1774
rect 877 -1735 881 -1731
rect 894 -1735 898 -1731
rect 628 -1848 632 -1844
rect 645 -1848 649 -1844
rect 1209 -1738 1213 -1734
rect 1226 -1738 1230 -1734
rect 2105 -1747 2109 -1743
rect 2127 -1747 2131 -1743
rect 2137 -1747 2141 -1743
rect 2159 -1747 2163 -1743
rect 1904 -1755 1908 -1751
rect 1926 -1755 1930 -1751
rect 1956 -1755 1960 -1751
rect 1978 -1755 1982 -1751
rect 2008 -1755 2012 -1751
rect 2030 -1755 2034 -1751
rect 2060 -1755 2064 -1751
rect 2082 -1755 2086 -1751
rect 1587 -1761 1591 -1757
rect 1604 -1761 1608 -1757
rect 1543 -1791 1547 -1787
rect 1543 -1808 1547 -1804
rect 1543 -1842 1547 -1838
rect 1543 -1859 1547 -1855
rect 554 -2027 558 -2023
rect 571 -2027 575 -2023
rect 581 -2027 585 -2023
rect 598 -2027 602 -2023
rect -275 -2108 -271 -2104
rect -253 -2108 -249 -2104
rect -243 -2108 -239 -2104
rect -221 -2108 -217 -2104
rect -476 -2116 -472 -2112
rect -454 -2116 -450 -2112
rect -424 -2116 -420 -2112
rect -402 -2116 -398 -2112
rect -372 -2116 -368 -2112
rect -350 -2116 -346 -2112
rect -320 -2116 -316 -2112
rect -298 -2116 -294 -2112
rect 616 -2097 620 -2093
rect 633 -2097 637 -2093
rect 206 -2327 210 -2323
rect 223 -2327 227 -2323
rect 1358 -2330 1362 -2326
rect 1375 -2330 1379 -2326
rect 162 -2357 166 -2353
rect 162 -2374 166 -2370
rect 693 -2337 697 -2333
rect 710 -2337 714 -2333
rect 720 -2337 724 -2333
rect 737 -2337 741 -2333
rect 162 -2408 166 -2404
rect 1028 -2389 1032 -2385
rect 1045 -2389 1049 -2385
rect 1055 -2389 1059 -2385
rect 1072 -2389 1076 -2385
rect 162 -2425 166 -2421
rect 123 -2471 127 -2467
rect 140 -2471 144 -2467
rect 150 -2471 154 -2467
rect 167 -2471 171 -2467
rect 755 -2407 759 -2403
rect 772 -2407 776 -2403
rect 2093 -2354 2097 -2350
rect 2110 -2354 2114 -2350
rect -266 -2537 -262 -2533
rect -244 -2537 -240 -2533
rect -234 -2537 -230 -2533
rect -212 -2537 -208 -2533
rect -467 -2545 -463 -2541
rect -445 -2545 -441 -2541
rect -415 -2545 -411 -2541
rect -393 -2545 -389 -2541
rect -363 -2545 -359 -2541
rect -341 -2545 -337 -2541
rect -311 -2545 -307 -2541
rect -289 -2545 -285 -2541
rect 1090 -2459 1094 -2455
rect 1107 -2459 1111 -2455
rect 185 -2541 189 -2537
rect 202 -2541 206 -2537
rect 2635 -2428 2639 -2424
rect 2657 -2428 2661 -2424
rect 2667 -2428 2671 -2424
rect 2689 -2428 2693 -2424
rect 2434 -2436 2438 -2432
rect 2456 -2436 2460 -2432
rect 2486 -2436 2490 -2432
rect 2508 -2436 2512 -2432
rect 2538 -2436 2542 -2432
rect 2560 -2436 2564 -2432
rect 2590 -2436 2594 -2432
rect 2612 -2436 2616 -2432
rect 1407 -2467 1411 -2463
rect 1424 -2467 1428 -2463
rect 2142 -2491 2146 -2487
rect 2159 -2491 2163 -2487
rect 694 -2620 698 -2616
rect 711 -2620 715 -2616
rect 721 -2620 725 -2616
rect 738 -2620 742 -2616
rect 1029 -2672 1033 -2668
rect 1046 -2672 1050 -2668
rect 1056 -2672 1060 -2668
rect 1073 -2672 1077 -2668
rect 756 -2690 760 -2686
rect 773 -2690 777 -2686
rect 1365 -2719 1369 -2715
rect 1382 -2719 1386 -2715
rect 1091 -2742 1095 -2738
rect 1108 -2742 1112 -2738
rect 690 -2891 694 -2887
rect 707 -2891 711 -2887
rect 717 -2891 721 -2887
rect 734 -2891 738 -2887
rect 1414 -2856 1418 -2852
rect 1431 -2856 1435 -2852
rect 1657 -2875 1661 -2871
rect 1674 -2875 1678 -2871
rect 752 -2961 756 -2957
rect 769 -2961 773 -2957
rect 1359 -3074 1363 -3070
rect 1376 -3074 1380 -3070
rect 1386 -3074 1390 -3070
rect 1403 -3074 1407 -3070
rect 1706 -3012 1710 -3008
rect 1723 -3012 1727 -3008
rect 678 -3140 682 -3136
rect 695 -3140 699 -3136
rect 705 -3140 709 -3136
rect 722 -3140 726 -3136
rect 1019 -3206 1023 -3202
rect 1036 -3206 1040 -3202
rect 1046 -3206 1050 -3202
rect 1063 -3206 1067 -3202
rect 740 -3210 744 -3206
rect 757 -3210 761 -3206
rect 1421 -3144 1425 -3140
rect 1438 -3144 1442 -3140
rect 1081 -3276 1085 -3272
rect 1098 -3276 1102 -3272
rect 695 -3407 699 -3403
rect 712 -3407 716 -3403
rect 722 -3407 726 -3403
rect 739 -3407 743 -3403
rect 757 -3477 761 -3473
rect 774 -3477 778 -3473
rect 683 -3656 687 -3652
rect 700 -3656 704 -3652
rect 710 -3656 714 -3652
rect 727 -3656 731 -3652
rect 745 -3726 749 -3722
rect 762 -3726 766 -3722
<< polysilicon >>
rect 1377 213 1379 217
rect 1409 213 1411 217
rect 1176 205 1178 209
rect 1228 205 1230 209
rect 1280 205 1282 209
rect 1332 205 1334 209
rect 1176 156 1178 165
rect 1228 156 1230 165
rect 1280 156 1282 165
rect 1332 156 1334 165
rect 1377 153 1379 173
rect 1409 153 1411 173
rect 1176 143 1178 147
rect 1228 143 1230 147
rect 1280 129 1282 138
rect 1332 129 1334 138
rect 1377 129 1379 133
rect 1409 129 1411 133
rect 1280 106 1282 109
rect 1332 106 1334 109
rect 1176 94 1178 103
rect 1228 94 1230 103
rect -254 87 -252 91
rect -222 87 -220 91
rect -455 79 -453 83
rect -403 79 -401 83
rect -351 79 -349 83
rect -299 79 -297 83
rect 1176 82 1178 90
rect 1228 82 1230 90
rect 1280 82 1282 90
rect 1332 82 1334 90
rect 1176 58 1178 62
rect 1228 58 1230 62
rect 1280 58 1282 62
rect 1332 58 1334 62
rect -455 30 -453 39
rect -403 30 -401 39
rect -351 30 -349 39
rect -299 30 -297 39
rect -254 27 -252 47
rect -222 27 -220 47
rect 515 27 597 29
rect 631 28 633 31
rect -455 17 -453 21
rect -403 17 -401 21
rect -351 3 -349 12
rect -299 3 -297 12
rect -254 3 -252 7
rect -222 3 -220 7
rect 595 5 597 27
rect 489 -3 492 -1
rect 512 -3 530 -1
rect 570 -3 573 -1
rect -351 -20 -349 -17
rect -299 -20 -297 -17
rect 595 -18 597 -15
rect -455 -32 -453 -23
rect -403 -32 -401 -23
rect 515 -25 597 -23
rect 595 -28 597 -25
rect -455 -44 -453 -36
rect -403 -44 -401 -36
rect -351 -44 -349 -36
rect -299 -44 -297 -36
rect 631 -30 633 -12
rect 595 -51 597 -48
rect 489 -54 492 -52
rect 512 -54 530 -52
rect 570 -54 573 -52
rect 631 -53 633 -50
rect -455 -68 -453 -64
rect -403 -68 -401 -64
rect -351 -68 -349 -64
rect -299 -68 -297 -64
rect 725 -146 727 -143
rect 143 -164 225 -162
rect 259 -163 261 -160
rect 223 -186 225 -164
rect 117 -194 120 -192
rect 140 -194 158 -192
rect 198 -194 201 -192
rect 480 -179 482 -176
rect 507 -179 509 -176
rect 223 -209 225 -206
rect 143 -216 225 -214
rect 223 -219 225 -216
rect 259 -221 261 -203
rect 223 -242 225 -239
rect 117 -245 120 -243
rect 140 -245 158 -243
rect 198 -245 201 -243
rect 259 -244 261 -241
rect 480 -247 482 -219
rect 507 -231 509 -219
rect 507 -233 517 -231
rect 480 -249 501 -247
rect 499 -253 501 -249
rect 499 -297 501 -293
rect -221 -308 -219 -304
rect -189 -308 -187 -304
rect 176 -307 178 -304
rect 203 -307 205 -304
rect -422 -316 -420 -312
rect -370 -316 -368 -312
rect -318 -316 -316 -312
rect -266 -316 -264 -312
rect 515 -310 517 -233
rect 725 -232 727 -226
rect 725 -234 745 -232
rect 725 -246 727 -243
rect 542 -249 544 -246
rect 542 -307 544 -289
rect 499 -312 517 -310
rect 499 -318 501 -312
rect -422 -365 -420 -356
rect -370 -365 -368 -356
rect -318 -365 -316 -356
rect -266 -365 -264 -356
rect -221 -368 -219 -348
rect -189 -368 -187 -348
rect -422 -378 -420 -374
rect -370 -378 -368 -374
rect -318 -392 -316 -383
rect -266 -392 -264 -383
rect 176 -375 178 -347
rect 203 -359 205 -347
rect 542 -330 544 -327
rect 725 -332 727 -326
rect 710 -334 727 -332
rect 710 -351 712 -334
rect 743 -351 745 -234
rect 1655 -250 1657 -246
rect 1687 -250 1689 -246
rect 1454 -258 1456 -254
rect 1506 -258 1508 -254
rect 1558 -258 1560 -254
rect 1610 -258 1612 -254
rect 774 -283 776 -280
rect 1454 -307 1456 -298
rect 1506 -307 1508 -298
rect 1558 -307 1560 -298
rect 1610 -307 1612 -298
rect 1655 -310 1657 -290
rect 1687 -310 1689 -290
rect 1454 -320 1456 -316
rect 1506 -320 1508 -316
rect 774 -341 776 -323
rect 203 -361 213 -359
rect 499 -361 501 -358
rect 176 -377 197 -375
rect 195 -381 197 -377
rect -221 -392 -219 -388
rect -189 -392 -187 -388
rect -318 -415 -316 -412
rect -266 -415 -264 -412
rect -422 -427 -420 -418
rect -370 -427 -368 -418
rect 195 -425 197 -421
rect -422 -439 -420 -431
rect -370 -439 -368 -431
rect -318 -439 -316 -431
rect -266 -439 -264 -431
rect 211 -438 213 -361
rect 1011 -360 1093 -358
rect 1127 -359 1129 -356
rect 774 -364 776 -361
rect 710 -374 712 -371
rect 743 -374 745 -371
rect 238 -377 240 -374
rect 1091 -382 1093 -360
rect 985 -390 988 -388
rect 1008 -390 1026 -388
rect 1066 -390 1069 -388
rect 1558 -334 1560 -325
rect 1610 -334 1612 -325
rect 1655 -334 1657 -330
rect 1687 -334 1689 -330
rect 1558 -357 1560 -354
rect 1610 -357 1612 -354
rect 1454 -369 1456 -360
rect 1506 -369 1508 -360
rect 1454 -381 1456 -373
rect 1506 -381 1508 -373
rect 1558 -381 1560 -373
rect 1610 -381 1612 -373
rect 1091 -405 1093 -402
rect 1011 -412 1093 -410
rect 1091 -415 1093 -412
rect 238 -435 240 -417
rect 195 -440 213 -438
rect 195 -446 197 -440
rect -422 -463 -420 -459
rect -370 -463 -368 -459
rect -318 -463 -316 -459
rect -266 -463 -264 -459
rect 1127 -417 1129 -399
rect 1454 -405 1456 -401
rect 1506 -405 1508 -401
rect 1558 -405 1560 -401
rect 1610 -405 1612 -401
rect 1091 -438 1093 -435
rect 985 -441 988 -439
rect 1008 -441 1026 -439
rect 1066 -441 1069 -439
rect 1127 -440 1129 -437
rect 238 -458 240 -455
rect 195 -489 197 -486
rect 1206 -627 1208 -624
rect 980 -635 982 -632
rect 581 -668 583 -665
rect 608 -668 610 -665
rect -330 -687 -328 -683
rect -298 -687 -296 -683
rect -531 -695 -529 -691
rect -479 -695 -477 -691
rect -427 -695 -425 -691
rect -375 -695 -373 -691
rect -531 -744 -529 -735
rect -479 -744 -477 -735
rect -427 -744 -425 -735
rect -375 -744 -373 -735
rect -330 -747 -328 -727
rect -298 -747 -296 -727
rect 581 -736 583 -708
rect 608 -720 610 -708
rect 1206 -713 1208 -707
rect 1206 -715 1226 -713
rect 608 -722 618 -720
rect 581 -738 602 -736
rect 600 -742 602 -738
rect -531 -757 -529 -753
rect -479 -757 -477 -753
rect -427 -771 -425 -762
rect -375 -771 -373 -762
rect -330 -771 -328 -767
rect -298 -771 -296 -767
rect 600 -786 602 -782
rect -427 -794 -425 -791
rect -375 -794 -373 -791
rect -531 -806 -529 -797
rect -479 -806 -477 -797
rect 94 -800 176 -798
rect 210 -799 212 -796
rect 616 -799 618 -722
rect 980 -721 982 -715
rect 980 -723 1000 -721
rect 980 -735 982 -732
rect 643 -738 645 -735
rect 643 -796 645 -778
rect -531 -818 -529 -810
rect -479 -818 -477 -810
rect -427 -818 -425 -810
rect -375 -818 -373 -810
rect 174 -822 176 -800
rect 68 -830 71 -828
rect 91 -830 109 -828
rect 149 -830 152 -828
rect -531 -842 -529 -838
rect -479 -842 -477 -838
rect -427 -842 -425 -838
rect -375 -842 -373 -838
rect 600 -801 618 -799
rect 600 -807 602 -801
rect 174 -845 176 -842
rect 94 -852 176 -850
rect 174 -855 176 -852
rect 210 -857 212 -839
rect 643 -819 645 -816
rect 980 -821 982 -815
rect 965 -823 982 -821
rect 965 -840 967 -823
rect 998 -840 1000 -723
rect 1206 -727 1208 -724
rect 1029 -772 1031 -769
rect 1029 -830 1031 -812
rect 1206 -813 1208 -807
rect 1191 -815 1208 -813
rect 600 -850 602 -847
rect 174 -878 176 -875
rect 1191 -832 1193 -815
rect 1224 -832 1226 -715
rect 1255 -764 1257 -761
rect 1255 -822 1257 -804
rect 1365 -805 1447 -803
rect 1481 -804 1483 -801
rect 1029 -853 1031 -850
rect 1445 -827 1447 -805
rect 1339 -835 1342 -833
rect 1362 -835 1380 -833
rect 1420 -835 1423 -833
rect 1255 -845 1257 -842
rect 1966 -805 1968 -801
rect 1998 -805 2000 -801
rect 1765 -813 1767 -809
rect 1817 -813 1819 -809
rect 1869 -813 1871 -809
rect 1921 -813 1923 -809
rect 1191 -855 1193 -852
rect 1224 -855 1226 -852
rect 1445 -850 1447 -847
rect 1365 -857 1447 -855
rect 965 -863 967 -860
rect 998 -863 1000 -860
rect 1445 -860 1447 -857
rect 68 -881 71 -879
rect 91 -881 109 -879
rect 149 -881 152 -879
rect 210 -880 212 -877
rect 1481 -862 1483 -844
rect 1765 -862 1767 -853
rect 1817 -862 1819 -853
rect 1869 -862 1871 -853
rect 1921 -862 1923 -853
rect 1445 -883 1447 -880
rect 1966 -865 1968 -845
rect 1998 -865 2000 -845
rect 1765 -875 1767 -871
rect 1817 -875 1819 -871
rect 1339 -886 1342 -884
rect 1362 -886 1380 -884
rect 1420 -886 1423 -884
rect 1481 -885 1483 -882
rect 504 -913 506 -910
rect 531 -913 533 -910
rect 722 -913 724 -910
rect 749 -913 751 -910
rect 127 -943 129 -940
rect 154 -943 156 -940
rect 1869 -889 1871 -880
rect 1921 -889 1923 -880
rect 1966 -889 1968 -885
rect 1998 -889 2000 -885
rect 1869 -912 1871 -909
rect 1921 -912 1923 -909
rect 1765 -924 1767 -915
rect 1817 -924 1819 -915
rect 1765 -936 1767 -928
rect 1817 -936 1819 -928
rect 1869 -936 1871 -928
rect 1921 -936 1923 -928
rect 504 -981 506 -953
rect 531 -965 533 -953
rect 531 -967 541 -965
rect 504 -983 525 -981
rect 127 -1011 129 -983
rect 154 -995 156 -983
rect 523 -987 525 -983
rect 154 -997 164 -995
rect 127 -1013 148 -1011
rect 146 -1017 148 -1013
rect -254 -1040 -252 -1036
rect -222 -1040 -220 -1036
rect -455 -1048 -453 -1044
rect -403 -1048 -401 -1044
rect -351 -1048 -349 -1044
rect -299 -1048 -297 -1044
rect 146 -1061 148 -1057
rect 162 -1074 164 -997
rect 189 -1013 191 -1010
rect 523 -1031 525 -1027
rect 539 -1044 541 -967
rect 566 -983 568 -980
rect 722 -981 724 -953
rect 749 -965 751 -953
rect 1765 -960 1767 -956
rect 1817 -960 1819 -956
rect 1869 -960 1871 -956
rect 1921 -960 1923 -956
rect 749 -967 759 -965
rect 722 -983 743 -981
rect 741 -987 743 -983
rect 566 -1041 568 -1023
rect 741 -1031 743 -1027
rect 523 -1046 541 -1044
rect 523 -1052 525 -1046
rect 189 -1071 191 -1053
rect 146 -1076 164 -1074
rect -455 -1097 -453 -1088
rect -403 -1097 -401 -1088
rect -351 -1097 -349 -1088
rect -299 -1097 -297 -1088
rect -254 -1100 -252 -1080
rect -222 -1100 -220 -1080
rect 146 -1082 148 -1076
rect -455 -1110 -453 -1106
rect -403 -1110 -401 -1106
rect -351 -1124 -349 -1115
rect -299 -1124 -297 -1115
rect -254 -1124 -252 -1120
rect -222 -1124 -220 -1120
rect 189 -1094 191 -1091
rect 757 -1044 759 -967
rect 784 -983 786 -980
rect 784 -1041 786 -1023
rect 741 -1046 759 -1044
rect 741 -1052 743 -1046
rect 566 -1064 568 -1061
rect 784 -1064 786 -1061
rect 523 -1095 525 -1092
rect 741 -1095 743 -1092
rect 146 -1125 148 -1122
rect -351 -1147 -349 -1144
rect -299 -1147 -297 -1144
rect -455 -1159 -453 -1150
rect -403 -1159 -401 -1150
rect -455 -1171 -453 -1163
rect -403 -1171 -401 -1163
rect -351 -1171 -349 -1163
rect -299 -1171 -297 -1163
rect -455 -1195 -453 -1191
rect -403 -1195 -401 -1191
rect -351 -1195 -349 -1191
rect -299 -1195 -297 -1191
rect 579 -1231 581 -1228
rect 606 -1231 608 -1228
rect 579 -1299 581 -1271
rect 606 -1283 608 -1271
rect 606 -1285 616 -1283
rect 579 -1301 600 -1299
rect 598 -1305 600 -1301
rect 598 -1349 600 -1345
rect 614 -1362 616 -1285
rect 641 -1301 643 -1298
rect 1159 -1308 1161 -1305
rect 641 -1359 643 -1341
rect -263 -1368 -261 -1364
rect -231 -1368 -229 -1364
rect 598 -1364 616 -1362
rect -464 -1376 -462 -1372
rect -412 -1376 -410 -1372
rect -360 -1376 -358 -1372
rect -308 -1376 -306 -1372
rect 598 -1370 600 -1364
rect -464 -1425 -462 -1416
rect -412 -1425 -410 -1416
rect -360 -1425 -358 -1416
rect -308 -1425 -306 -1416
rect -263 -1428 -261 -1408
rect -231 -1428 -229 -1408
rect 641 -1382 643 -1379
rect 1159 -1394 1161 -1388
rect 1159 -1396 1179 -1394
rect 1159 -1408 1161 -1405
rect 598 -1413 600 -1410
rect -464 -1438 -462 -1434
rect -412 -1438 -410 -1434
rect -360 -1452 -358 -1443
rect -308 -1452 -306 -1443
rect -263 -1452 -261 -1448
rect -231 -1452 -229 -1448
rect 103 -1460 185 -1458
rect 219 -1459 221 -1456
rect -360 -1475 -358 -1472
rect -308 -1475 -306 -1472
rect -464 -1487 -462 -1478
rect -412 -1487 -410 -1478
rect 183 -1482 185 -1460
rect 77 -1490 80 -1488
rect 100 -1490 118 -1488
rect 158 -1490 161 -1488
rect -464 -1499 -462 -1491
rect -412 -1499 -410 -1491
rect -360 -1499 -358 -1491
rect -308 -1499 -306 -1491
rect 816 -1461 818 -1458
rect 843 -1461 845 -1458
rect 183 -1505 185 -1502
rect 103 -1512 185 -1510
rect 183 -1515 185 -1512
rect -464 -1523 -462 -1519
rect -412 -1523 -410 -1519
rect -360 -1523 -358 -1519
rect -308 -1523 -306 -1519
rect 219 -1517 221 -1499
rect 1159 -1494 1161 -1488
rect 1144 -1496 1161 -1494
rect 580 -1514 582 -1511
rect 607 -1514 609 -1511
rect 183 -1538 185 -1535
rect 77 -1541 80 -1539
rect 100 -1541 118 -1539
rect 158 -1541 161 -1539
rect 219 -1540 221 -1537
rect 816 -1529 818 -1501
rect 843 -1513 845 -1501
rect 1144 -1513 1146 -1496
rect 1177 -1513 1179 -1396
rect 1208 -1445 1210 -1442
rect 1319 -1472 1321 -1469
rect 1208 -1503 1210 -1485
rect 843 -1515 853 -1513
rect 816 -1531 837 -1529
rect 835 -1535 837 -1531
rect 580 -1582 582 -1554
rect 607 -1566 609 -1554
rect 607 -1568 617 -1566
rect 580 -1584 601 -1582
rect 599 -1588 601 -1584
rect 136 -1603 138 -1600
rect 163 -1603 165 -1600
rect 599 -1632 601 -1628
rect 136 -1671 138 -1643
rect 163 -1655 165 -1643
rect 615 -1645 617 -1568
rect 835 -1579 837 -1575
rect 642 -1584 644 -1581
rect 851 -1592 853 -1515
rect 878 -1531 880 -1528
rect 1208 -1526 1210 -1523
rect 1144 -1536 1146 -1533
rect 1177 -1536 1179 -1533
rect 1319 -1558 1321 -1552
rect 1319 -1560 1339 -1558
rect 878 -1589 880 -1571
rect 1319 -1572 1321 -1569
rect 835 -1594 853 -1592
rect 835 -1600 837 -1594
rect 642 -1642 644 -1624
rect 1170 -1608 1172 -1605
rect 878 -1612 880 -1609
rect 599 -1647 617 -1645
rect 599 -1653 601 -1647
rect 163 -1657 173 -1655
rect 136 -1673 157 -1671
rect 155 -1677 157 -1673
rect 155 -1721 157 -1717
rect 171 -1734 173 -1657
rect 198 -1673 200 -1670
rect 835 -1643 837 -1640
rect 642 -1665 644 -1662
rect 825 -1672 827 -1669
rect 852 -1672 854 -1669
rect 599 -1696 601 -1693
rect 1319 -1658 1321 -1652
rect 1304 -1660 1321 -1658
rect 1304 -1677 1306 -1660
rect 1337 -1677 1339 -1560
rect 1368 -1609 1370 -1606
rect 1368 -1667 1370 -1649
rect 1170 -1694 1172 -1688
rect 1170 -1696 1190 -1694
rect 1170 -1708 1172 -1705
rect 198 -1731 200 -1713
rect 155 -1736 173 -1734
rect 155 -1742 157 -1736
rect -279 -1746 -277 -1742
rect -247 -1746 -245 -1742
rect -480 -1754 -478 -1750
rect -428 -1754 -426 -1750
rect -376 -1754 -374 -1750
rect -324 -1754 -322 -1750
rect 825 -1740 827 -1712
rect 852 -1724 854 -1712
rect 852 -1726 862 -1724
rect 825 -1742 846 -1740
rect 844 -1746 846 -1742
rect 198 -1754 200 -1751
rect 155 -1785 157 -1782
rect 576 -1785 578 -1782
rect 603 -1785 605 -1782
rect -480 -1803 -478 -1794
rect -428 -1803 -426 -1794
rect -376 -1803 -374 -1794
rect -324 -1803 -322 -1794
rect -279 -1806 -277 -1786
rect -247 -1806 -245 -1786
rect -480 -1816 -478 -1812
rect -428 -1816 -426 -1812
rect -376 -1830 -374 -1821
rect -324 -1830 -322 -1821
rect 844 -1790 846 -1786
rect 860 -1803 862 -1726
rect 887 -1742 889 -1739
rect 887 -1800 889 -1782
rect 1170 -1794 1172 -1788
rect 1155 -1796 1172 -1794
rect 844 -1805 862 -1803
rect 844 -1811 846 -1805
rect -279 -1830 -277 -1826
rect -247 -1830 -245 -1826
rect -376 -1853 -374 -1850
rect -324 -1853 -322 -1850
rect 576 -1853 578 -1825
rect 603 -1837 605 -1825
rect 603 -1839 613 -1837
rect 576 -1855 597 -1853
rect -480 -1865 -478 -1856
rect -428 -1865 -426 -1856
rect 595 -1859 597 -1855
rect -480 -1877 -478 -1869
rect -428 -1877 -426 -1869
rect -376 -1877 -374 -1869
rect -324 -1877 -322 -1869
rect -480 -1901 -478 -1897
rect -428 -1901 -426 -1897
rect -376 -1901 -374 -1897
rect -324 -1901 -322 -1897
rect 595 -1903 597 -1899
rect 611 -1916 613 -1839
rect 1155 -1813 1157 -1796
rect 1188 -1813 1190 -1696
rect 1368 -1690 1370 -1687
rect 1304 -1700 1306 -1697
rect 1337 -1700 1339 -1697
rect 1219 -1745 1221 -1742
rect 2117 -1755 2119 -1751
rect 2149 -1755 2151 -1751
rect 1916 -1763 1918 -1759
rect 1968 -1763 1970 -1759
rect 2020 -1763 2022 -1759
rect 2072 -1763 2074 -1759
rect 1481 -1769 1563 -1767
rect 1597 -1768 1599 -1765
rect 1219 -1803 1221 -1785
rect 1561 -1791 1563 -1769
rect 1455 -1799 1458 -1797
rect 1478 -1799 1496 -1797
rect 1536 -1799 1539 -1797
rect 887 -1823 889 -1820
rect 1561 -1814 1563 -1811
rect 1481 -1821 1563 -1819
rect 1219 -1826 1221 -1823
rect 1561 -1824 1563 -1821
rect 1155 -1836 1157 -1833
rect 1188 -1836 1190 -1833
rect 1597 -1826 1599 -1808
rect 1916 -1812 1918 -1803
rect 1968 -1812 1970 -1803
rect 2020 -1812 2022 -1803
rect 2072 -1812 2074 -1803
rect 2117 -1815 2119 -1795
rect 2149 -1815 2151 -1795
rect 1916 -1825 1918 -1821
rect 1968 -1825 1970 -1821
rect 1561 -1847 1563 -1844
rect 1455 -1850 1458 -1848
rect 1478 -1850 1496 -1848
rect 1536 -1850 1539 -1848
rect 1597 -1849 1599 -1846
rect 638 -1855 640 -1852
rect 844 -1854 846 -1851
rect 2020 -1839 2022 -1830
rect 2072 -1839 2074 -1830
rect 2117 -1839 2119 -1835
rect 2149 -1839 2151 -1835
rect 2020 -1862 2022 -1859
rect 2072 -1862 2074 -1859
rect 1916 -1874 1918 -1865
rect 1968 -1874 1970 -1865
rect 1916 -1886 1918 -1878
rect 1968 -1886 1970 -1878
rect 2020 -1886 2022 -1878
rect 2072 -1886 2074 -1878
rect 638 -1913 640 -1895
rect 1916 -1910 1918 -1906
rect 1968 -1910 1970 -1906
rect 2020 -1910 2022 -1906
rect 2072 -1910 2074 -1906
rect 595 -1918 613 -1916
rect 595 -1924 597 -1918
rect 638 -1936 640 -1933
rect 595 -1967 597 -1964
rect 564 -2034 566 -2031
rect 591 -2034 593 -2031
rect 564 -2102 566 -2074
rect 591 -2086 593 -2074
rect 591 -2088 601 -2086
rect 564 -2104 585 -2102
rect 583 -2108 585 -2104
rect -263 -2116 -261 -2112
rect -231 -2116 -229 -2112
rect -464 -2124 -462 -2120
rect -412 -2124 -410 -2120
rect -360 -2124 -358 -2120
rect -308 -2124 -306 -2120
rect 583 -2152 585 -2148
rect -464 -2173 -462 -2164
rect -412 -2173 -410 -2164
rect -360 -2173 -358 -2164
rect -308 -2173 -306 -2164
rect -263 -2176 -261 -2156
rect -231 -2176 -229 -2156
rect 599 -2165 601 -2088
rect 626 -2104 628 -2101
rect 626 -2162 628 -2144
rect 583 -2167 601 -2165
rect 583 -2173 585 -2167
rect -464 -2186 -462 -2182
rect -412 -2186 -410 -2182
rect -360 -2200 -358 -2191
rect -308 -2200 -306 -2191
rect -263 -2200 -261 -2196
rect -231 -2200 -229 -2196
rect 626 -2185 628 -2182
rect 583 -2216 585 -2213
rect -360 -2223 -358 -2220
rect -308 -2223 -306 -2220
rect -464 -2235 -462 -2226
rect -412 -2235 -410 -2226
rect -464 -2247 -462 -2239
rect -412 -2247 -410 -2239
rect -360 -2247 -358 -2239
rect -308 -2247 -306 -2239
rect -464 -2271 -462 -2267
rect -412 -2271 -410 -2267
rect -360 -2271 -358 -2267
rect -308 -2271 -306 -2267
rect 100 -2335 182 -2333
rect 216 -2334 218 -2331
rect 180 -2357 182 -2335
rect 74 -2365 77 -2363
rect 97 -2365 115 -2363
rect 155 -2365 158 -2363
rect 1368 -2337 1370 -2334
rect 703 -2344 705 -2341
rect 730 -2344 732 -2341
rect 180 -2380 182 -2377
rect 100 -2387 182 -2385
rect 180 -2390 182 -2387
rect 216 -2392 218 -2374
rect 180 -2413 182 -2410
rect 74 -2416 77 -2414
rect 97 -2416 115 -2414
rect 155 -2416 158 -2414
rect 216 -2415 218 -2412
rect 703 -2412 705 -2384
rect 730 -2396 732 -2384
rect 1038 -2396 1040 -2393
rect 1065 -2396 1067 -2393
rect 730 -2398 740 -2396
rect 703 -2414 724 -2412
rect 722 -2418 724 -2414
rect 722 -2462 724 -2458
rect 738 -2475 740 -2398
rect 765 -2414 767 -2411
rect 2103 -2361 2105 -2358
rect 1368 -2423 1370 -2417
rect 1368 -2425 1388 -2423
rect 765 -2472 767 -2454
rect 1038 -2464 1040 -2436
rect 1065 -2448 1067 -2436
rect 1368 -2437 1370 -2434
rect 1065 -2450 1075 -2448
rect 1038 -2466 1059 -2464
rect 1057 -2470 1059 -2466
rect 133 -2478 135 -2475
rect 160 -2478 162 -2475
rect 722 -2477 740 -2475
rect 722 -2483 724 -2477
rect -254 -2545 -252 -2541
rect -222 -2545 -220 -2541
rect -455 -2553 -453 -2549
rect -403 -2553 -401 -2549
rect -351 -2553 -349 -2549
rect -299 -2553 -297 -2549
rect 133 -2546 135 -2518
rect 160 -2530 162 -2518
rect 765 -2495 767 -2492
rect 1057 -2514 1059 -2510
rect 722 -2526 724 -2523
rect 1073 -2527 1075 -2450
rect 1100 -2466 1102 -2463
rect 1100 -2524 1102 -2506
rect 1368 -2523 1370 -2517
rect 160 -2532 170 -2530
rect 133 -2548 154 -2546
rect 152 -2552 154 -2548
rect -455 -2602 -453 -2593
rect -403 -2602 -401 -2593
rect -351 -2602 -349 -2593
rect -299 -2602 -297 -2593
rect -254 -2605 -252 -2585
rect -222 -2605 -220 -2585
rect 152 -2596 154 -2592
rect -455 -2615 -453 -2611
rect -403 -2615 -401 -2611
rect -351 -2629 -349 -2620
rect -299 -2629 -297 -2620
rect 168 -2609 170 -2532
rect 1057 -2529 1075 -2527
rect 1057 -2535 1059 -2529
rect 195 -2548 197 -2545
rect 1353 -2525 1370 -2523
rect 1353 -2542 1355 -2525
rect 1386 -2542 1388 -2425
rect 2647 -2436 2649 -2432
rect 2679 -2436 2681 -2432
rect 2103 -2447 2105 -2441
rect 2446 -2444 2448 -2440
rect 2498 -2444 2500 -2440
rect 2550 -2444 2552 -2440
rect 2602 -2444 2604 -2440
rect 2103 -2449 2123 -2447
rect 2103 -2461 2105 -2458
rect 1417 -2474 1419 -2471
rect 1417 -2532 1419 -2514
rect 1100 -2547 1102 -2544
rect 2103 -2547 2105 -2541
rect 2088 -2549 2105 -2547
rect 1417 -2555 1419 -2552
rect 1353 -2565 1355 -2562
rect 1386 -2565 1388 -2562
rect 2088 -2566 2090 -2549
rect 2121 -2566 2123 -2449
rect 2446 -2493 2448 -2484
rect 2498 -2493 2500 -2484
rect 2550 -2493 2552 -2484
rect 2602 -2493 2604 -2484
rect 2152 -2498 2154 -2495
rect 2647 -2496 2649 -2476
rect 2679 -2496 2681 -2476
rect 2446 -2506 2448 -2502
rect 2498 -2506 2500 -2502
rect 2152 -2556 2154 -2538
rect 2550 -2520 2552 -2511
rect 2602 -2520 2604 -2511
rect 2647 -2520 2649 -2516
rect 2679 -2520 2681 -2516
rect 2550 -2543 2552 -2540
rect 2602 -2543 2604 -2540
rect 2446 -2555 2448 -2546
rect 2498 -2555 2500 -2546
rect 1057 -2578 1059 -2575
rect 2446 -2567 2448 -2559
rect 2498 -2567 2500 -2559
rect 2550 -2567 2552 -2559
rect 2602 -2567 2604 -2559
rect 2152 -2579 2154 -2576
rect 195 -2606 197 -2588
rect 2088 -2589 2090 -2586
rect 2121 -2589 2123 -2586
rect 2446 -2591 2448 -2587
rect 2498 -2591 2500 -2587
rect 2550 -2591 2552 -2587
rect 2602 -2591 2604 -2587
rect 152 -2611 170 -2609
rect 152 -2617 154 -2611
rect -254 -2629 -252 -2625
rect -222 -2629 -220 -2625
rect -351 -2652 -349 -2649
rect -299 -2652 -297 -2649
rect -455 -2664 -453 -2655
rect -403 -2664 -401 -2655
rect 195 -2629 197 -2626
rect 704 -2627 706 -2624
rect 731 -2627 733 -2624
rect 152 -2660 154 -2657
rect -455 -2676 -453 -2668
rect -403 -2676 -401 -2668
rect -351 -2676 -349 -2668
rect -299 -2676 -297 -2668
rect -455 -2700 -453 -2696
rect -403 -2700 -401 -2696
rect -351 -2700 -349 -2696
rect -299 -2700 -297 -2696
rect 704 -2695 706 -2667
rect 731 -2679 733 -2667
rect 1039 -2679 1041 -2676
rect 1066 -2679 1068 -2676
rect 731 -2681 741 -2679
rect 704 -2697 725 -2695
rect 723 -2701 725 -2697
rect 723 -2745 725 -2741
rect 739 -2758 741 -2681
rect 766 -2697 768 -2694
rect 766 -2755 768 -2737
rect 1039 -2747 1041 -2719
rect 1066 -2731 1068 -2719
rect 1375 -2726 1377 -2723
rect 1066 -2733 1076 -2731
rect 1039 -2749 1060 -2747
rect 1058 -2753 1060 -2749
rect 723 -2760 741 -2758
rect 723 -2766 725 -2760
rect 766 -2778 768 -2775
rect 1058 -2797 1060 -2793
rect 723 -2809 725 -2806
rect 1074 -2810 1076 -2733
rect 1101 -2749 1103 -2746
rect 1101 -2807 1103 -2789
rect 1058 -2812 1076 -2810
rect 1058 -2818 1060 -2812
rect 1375 -2812 1377 -2806
rect 1375 -2814 1395 -2812
rect 1375 -2826 1377 -2823
rect 1101 -2830 1103 -2827
rect 1058 -2861 1060 -2858
rect 700 -2898 702 -2895
rect 727 -2898 729 -2895
rect 1375 -2912 1377 -2906
rect 1360 -2914 1377 -2912
rect 1360 -2931 1362 -2914
rect 1393 -2931 1395 -2814
rect 1424 -2863 1426 -2860
rect 1667 -2882 1669 -2879
rect 1424 -2921 1426 -2903
rect 700 -2966 702 -2938
rect 727 -2950 729 -2938
rect 727 -2952 737 -2950
rect 1424 -2944 1426 -2941
rect 700 -2968 721 -2966
rect 719 -2972 721 -2968
rect 719 -3016 721 -3012
rect 735 -3029 737 -2952
rect 1360 -2954 1362 -2951
rect 1393 -2954 1395 -2951
rect 762 -2968 764 -2965
rect 1667 -2968 1669 -2962
rect 1667 -2970 1687 -2968
rect 1667 -2982 1669 -2979
rect 762 -3026 764 -3008
rect 719 -3031 737 -3029
rect 719 -3037 721 -3031
rect 762 -3049 764 -3046
rect 1667 -3068 1669 -3062
rect 1652 -3070 1669 -3068
rect 719 -3080 721 -3077
rect 1369 -3081 1371 -3078
rect 1396 -3081 1398 -3078
rect 1652 -3087 1654 -3070
rect 1685 -3087 1687 -2970
rect 1716 -3019 1718 -3016
rect 1716 -3077 1718 -3059
rect 1716 -3100 1718 -3097
rect 1652 -3110 1654 -3107
rect 1685 -3110 1687 -3107
rect 688 -3147 690 -3144
rect 715 -3147 717 -3144
rect 1369 -3149 1371 -3121
rect 1396 -3133 1398 -3121
rect 1396 -3135 1406 -3133
rect 1369 -3151 1390 -3149
rect 1388 -3155 1390 -3151
rect 688 -3215 690 -3187
rect 715 -3199 717 -3187
rect 1388 -3199 1390 -3195
rect 715 -3201 725 -3199
rect 688 -3217 709 -3215
rect 707 -3221 709 -3217
rect 707 -3265 709 -3261
rect 723 -3278 725 -3201
rect 1029 -3213 1031 -3210
rect 1056 -3213 1058 -3210
rect 1404 -3212 1406 -3135
rect 1431 -3151 1433 -3148
rect 1431 -3209 1433 -3191
rect 750 -3217 752 -3214
rect 1388 -3214 1406 -3212
rect 1388 -3220 1390 -3214
rect 750 -3275 752 -3257
rect 707 -3280 725 -3278
rect 707 -3286 709 -3280
rect 1029 -3281 1031 -3253
rect 1056 -3265 1058 -3253
rect 1431 -3232 1433 -3229
rect 1388 -3263 1390 -3260
rect 1056 -3267 1066 -3265
rect 1029 -3283 1050 -3281
rect 1048 -3287 1050 -3283
rect 750 -3298 752 -3295
rect 707 -3329 709 -3326
rect 1048 -3331 1050 -3327
rect 1064 -3344 1066 -3267
rect 1091 -3283 1093 -3280
rect 1091 -3341 1093 -3323
rect 1048 -3346 1066 -3344
rect 1048 -3352 1050 -3346
rect 1091 -3364 1093 -3361
rect 1048 -3395 1050 -3392
rect 705 -3414 707 -3411
rect 732 -3414 734 -3411
rect 705 -3482 707 -3454
rect 732 -3466 734 -3454
rect 732 -3468 742 -3466
rect 705 -3484 726 -3482
rect 724 -3488 726 -3484
rect 724 -3532 726 -3528
rect 740 -3545 742 -3468
rect 767 -3484 769 -3481
rect 767 -3542 769 -3524
rect 724 -3547 742 -3545
rect 724 -3553 726 -3547
rect 767 -3565 769 -3562
rect 724 -3596 726 -3593
rect 693 -3663 695 -3660
rect 720 -3663 722 -3660
rect 693 -3731 695 -3703
rect 720 -3715 722 -3703
rect 720 -3717 730 -3715
rect 693 -3733 714 -3731
rect 712 -3737 714 -3733
rect 712 -3781 714 -3777
rect 728 -3794 730 -3717
rect 755 -3733 757 -3730
rect 755 -3791 757 -3773
rect 712 -3796 730 -3794
rect 712 -3802 714 -3796
rect 755 -3814 757 -3811
rect 712 -3845 714 -3842
<< polycontact >>
rect 1171 156 1176 161
rect 1223 156 1228 161
rect 1275 156 1280 161
rect 1327 156 1332 161
rect 1372 156 1377 161
rect 1404 156 1409 161
rect 1275 133 1280 138
rect 1327 133 1332 138
rect 1171 94 1176 99
rect 1223 94 1228 99
rect 1171 85 1176 90
rect 1223 85 1228 90
rect 1275 85 1280 90
rect 1327 85 1332 90
rect -460 30 -455 35
rect -408 30 -403 35
rect -356 30 -351 35
rect -304 30 -299 35
rect -259 30 -254 35
rect -227 30 -222 35
rect -356 7 -351 12
rect -304 7 -299 12
rect 515 22 520 27
rect 515 -1 520 4
rect 515 -23 520 -18
rect -460 -32 -455 -27
rect -408 -32 -403 -27
rect 626 -27 631 -22
rect -460 -41 -455 -36
rect -408 -41 -403 -36
rect -356 -41 -351 -36
rect -304 -41 -299 -36
rect 515 -52 520 -47
rect 143 -169 148 -164
rect 143 -192 148 -187
rect 143 -214 148 -209
rect 254 -218 259 -213
rect 143 -243 148 -238
rect 475 -249 480 -244
rect 720 -234 725 -229
rect 537 -304 542 -299
rect 494 -315 499 -310
rect -427 -365 -422 -360
rect -375 -365 -370 -360
rect -323 -365 -318 -360
rect -271 -365 -266 -360
rect -226 -365 -221 -360
rect -194 -365 -189 -360
rect -323 -388 -318 -383
rect -271 -388 -266 -383
rect 171 -377 176 -372
rect 705 -337 710 -332
rect 1449 -307 1454 -302
rect 1501 -307 1506 -302
rect 1553 -307 1558 -302
rect 1605 -307 1610 -302
rect 1650 -307 1655 -302
rect 1682 -307 1687 -302
rect 769 -338 774 -333
rect -427 -427 -422 -422
rect -375 -427 -370 -422
rect -427 -436 -422 -431
rect -375 -436 -370 -431
rect -323 -436 -318 -431
rect -271 -436 -266 -431
rect 1011 -365 1016 -360
rect 1011 -388 1016 -383
rect 1553 -330 1558 -325
rect 1605 -330 1610 -325
rect 1449 -369 1454 -364
rect 1501 -369 1506 -364
rect 1449 -378 1454 -373
rect 1501 -378 1506 -373
rect 1553 -378 1558 -373
rect 1605 -378 1610 -373
rect 1011 -410 1016 -405
rect 1122 -414 1127 -409
rect 233 -432 238 -427
rect 190 -443 195 -438
rect 1011 -439 1016 -434
rect -536 -744 -531 -739
rect -484 -744 -479 -739
rect -432 -744 -427 -739
rect -380 -744 -375 -739
rect -335 -744 -330 -739
rect -303 -744 -298 -739
rect 576 -738 581 -733
rect 1201 -715 1206 -710
rect -432 -767 -427 -762
rect -380 -767 -375 -762
rect -536 -806 -531 -801
rect -484 -806 -479 -801
rect 975 -723 980 -718
rect 638 -793 643 -788
rect 94 -805 99 -800
rect -536 -815 -531 -810
rect -484 -815 -479 -810
rect -432 -815 -427 -810
rect -380 -815 -375 -810
rect 94 -828 99 -823
rect 595 -804 600 -799
rect 94 -850 99 -845
rect 205 -854 210 -849
rect 94 -879 99 -874
rect 960 -826 965 -821
rect 1024 -827 1029 -822
rect 1186 -818 1191 -813
rect 1250 -819 1255 -814
rect 1365 -810 1370 -805
rect 1365 -833 1370 -828
rect 1365 -855 1370 -850
rect 1476 -859 1481 -854
rect 1365 -884 1370 -879
rect 1760 -862 1765 -857
rect 1812 -862 1817 -857
rect 1864 -862 1869 -857
rect 1916 -862 1921 -857
rect 1961 -862 1966 -857
rect 1993 -862 1998 -857
rect 1864 -885 1869 -880
rect 1916 -885 1921 -880
rect 1760 -924 1765 -919
rect 1812 -924 1817 -919
rect 1760 -933 1765 -928
rect 1812 -933 1817 -928
rect 1864 -933 1869 -928
rect 1916 -933 1921 -928
rect 499 -983 504 -978
rect 122 -1013 127 -1008
rect 717 -983 722 -978
rect 561 -1038 566 -1033
rect 518 -1049 523 -1044
rect 184 -1068 189 -1063
rect 141 -1079 146 -1074
rect -460 -1097 -455 -1092
rect -408 -1097 -403 -1092
rect -356 -1097 -351 -1092
rect -304 -1097 -299 -1092
rect -259 -1097 -254 -1092
rect -227 -1097 -222 -1092
rect -356 -1120 -351 -1115
rect -304 -1120 -299 -1115
rect 779 -1038 784 -1033
rect 736 -1049 741 -1044
rect -460 -1159 -455 -1154
rect -408 -1159 -403 -1154
rect -460 -1168 -455 -1163
rect -408 -1168 -403 -1163
rect -356 -1168 -351 -1163
rect -304 -1168 -299 -1163
rect 574 -1301 579 -1296
rect 636 -1356 641 -1351
rect 593 -1367 598 -1362
rect -469 -1425 -464 -1420
rect -417 -1425 -412 -1420
rect -365 -1425 -360 -1420
rect -313 -1425 -308 -1420
rect -268 -1425 -263 -1420
rect -236 -1425 -231 -1420
rect 1154 -1396 1159 -1391
rect -365 -1448 -360 -1443
rect -313 -1448 -308 -1443
rect 103 -1465 108 -1460
rect -469 -1487 -464 -1482
rect -417 -1487 -412 -1482
rect 103 -1488 108 -1483
rect -469 -1496 -464 -1491
rect -417 -1496 -412 -1491
rect -365 -1496 -360 -1491
rect -313 -1496 -308 -1491
rect 103 -1510 108 -1505
rect 214 -1514 219 -1509
rect 103 -1539 108 -1534
rect 1139 -1499 1144 -1494
rect 811 -1531 816 -1526
rect 1203 -1500 1208 -1495
rect 575 -1584 580 -1579
rect 131 -1673 136 -1668
rect 1314 -1560 1319 -1555
rect 873 -1586 878 -1581
rect 830 -1597 835 -1592
rect 637 -1639 642 -1634
rect 594 -1650 599 -1645
rect 1299 -1663 1304 -1658
rect 1363 -1664 1368 -1659
rect 1165 -1696 1170 -1691
rect 193 -1728 198 -1723
rect 150 -1739 155 -1734
rect 820 -1742 825 -1737
rect -485 -1803 -480 -1798
rect -433 -1803 -428 -1798
rect -381 -1803 -376 -1798
rect -329 -1803 -324 -1798
rect -284 -1803 -279 -1798
rect -252 -1803 -247 -1798
rect -381 -1826 -376 -1821
rect -329 -1826 -324 -1821
rect 882 -1797 887 -1792
rect 1150 -1799 1155 -1794
rect 839 -1808 844 -1803
rect 571 -1855 576 -1850
rect -485 -1865 -480 -1860
rect -433 -1865 -428 -1860
rect -485 -1874 -480 -1869
rect -433 -1874 -428 -1869
rect -381 -1874 -376 -1869
rect -329 -1874 -324 -1869
rect 1481 -1774 1486 -1769
rect 1214 -1800 1219 -1795
rect 1481 -1797 1486 -1792
rect 1481 -1819 1486 -1814
rect 1592 -1823 1597 -1818
rect 1481 -1848 1486 -1843
rect 1911 -1812 1916 -1807
rect 1963 -1812 1968 -1807
rect 2015 -1812 2020 -1807
rect 2067 -1812 2072 -1807
rect 2112 -1812 2117 -1807
rect 2144 -1812 2149 -1807
rect 2015 -1835 2020 -1830
rect 2067 -1835 2072 -1830
rect 1911 -1874 1916 -1869
rect 1963 -1874 1968 -1869
rect 1911 -1883 1916 -1878
rect 1963 -1883 1968 -1878
rect 2015 -1883 2020 -1878
rect 2067 -1883 2072 -1878
rect 633 -1910 638 -1905
rect 590 -1921 595 -1916
rect 559 -2104 564 -2099
rect -469 -2173 -464 -2168
rect -417 -2173 -412 -2168
rect -365 -2173 -360 -2168
rect -313 -2173 -308 -2168
rect -268 -2173 -263 -2168
rect -236 -2173 -231 -2168
rect 621 -2159 626 -2154
rect 578 -2170 583 -2165
rect -365 -2196 -360 -2191
rect -313 -2196 -308 -2191
rect -469 -2235 -464 -2230
rect -417 -2235 -412 -2230
rect -469 -2244 -464 -2239
rect -417 -2244 -412 -2239
rect -365 -2244 -360 -2239
rect -313 -2244 -308 -2239
rect 100 -2340 105 -2335
rect 100 -2363 105 -2358
rect 100 -2385 105 -2380
rect 211 -2389 216 -2384
rect 100 -2414 105 -2409
rect 698 -2414 703 -2409
rect 1363 -2425 1368 -2420
rect 760 -2469 765 -2464
rect 1033 -2466 1038 -2461
rect 717 -2480 722 -2475
rect 128 -2548 133 -2543
rect 1095 -2521 1100 -2516
rect -460 -2602 -455 -2597
rect -408 -2602 -403 -2597
rect -356 -2602 -351 -2597
rect -304 -2602 -299 -2597
rect -259 -2602 -254 -2597
rect -227 -2602 -222 -2597
rect -356 -2625 -351 -2620
rect -304 -2625 -299 -2620
rect 1052 -2532 1057 -2527
rect 1348 -2528 1353 -2523
rect 2098 -2449 2103 -2444
rect 1412 -2529 1417 -2524
rect 2083 -2552 2088 -2547
rect 2441 -2493 2446 -2488
rect 2493 -2493 2498 -2488
rect 2545 -2493 2550 -2488
rect 2597 -2493 2602 -2488
rect 2642 -2493 2647 -2488
rect 2674 -2493 2679 -2488
rect 2147 -2553 2152 -2548
rect 2545 -2516 2550 -2511
rect 2597 -2516 2602 -2511
rect 2441 -2555 2446 -2550
rect 2493 -2555 2498 -2550
rect 2441 -2564 2446 -2559
rect 2493 -2564 2498 -2559
rect 2545 -2564 2550 -2559
rect 2597 -2564 2602 -2559
rect 190 -2603 195 -2598
rect 147 -2614 152 -2609
rect -460 -2664 -455 -2659
rect -408 -2664 -403 -2659
rect -460 -2673 -455 -2668
rect -408 -2673 -403 -2668
rect -356 -2673 -351 -2668
rect -304 -2673 -299 -2668
rect 699 -2697 704 -2692
rect 761 -2752 766 -2747
rect 1034 -2749 1039 -2744
rect 718 -2763 723 -2758
rect 1096 -2804 1101 -2799
rect 1053 -2815 1058 -2810
rect 1370 -2814 1375 -2809
rect 1355 -2917 1360 -2912
rect 1419 -2918 1424 -2913
rect 695 -2968 700 -2963
rect 1662 -2970 1667 -2965
rect 757 -3023 762 -3018
rect 714 -3034 719 -3029
rect 1647 -3073 1652 -3068
rect 1711 -3074 1716 -3069
rect 1364 -3151 1369 -3146
rect 683 -3217 688 -3212
rect 1426 -3206 1431 -3201
rect 1383 -3217 1388 -3212
rect 745 -3272 750 -3267
rect 702 -3283 707 -3278
rect 1024 -3283 1029 -3278
rect 1086 -3338 1091 -3333
rect 1043 -3349 1048 -3344
rect 700 -3484 705 -3479
rect 762 -3539 767 -3534
rect 719 -3550 724 -3545
rect 688 -3733 693 -3728
rect 750 -3788 755 -3783
rect 707 -3799 712 -3794
<< metal1 >>
rect 1362 225 1426 228
rect 1362 221 1365 225
rect 1369 221 1387 225
rect 1391 221 1397 225
rect 1401 221 1419 225
rect 1423 221 1426 225
rect 1161 217 1349 220
rect 1362 219 1426 221
rect 1161 213 1164 217
rect 1168 213 1186 217
rect 1190 213 1216 217
rect 1220 213 1238 217
rect 1242 213 1268 217
rect 1272 213 1290 217
rect 1294 213 1320 217
rect 1324 213 1342 217
rect 1346 213 1349 217
rect 1161 211 1349 213
rect 1372 213 1376 219
rect 1404 213 1408 219
rect 1171 205 1175 211
rect 1223 205 1227 211
rect 1275 205 1279 211
rect 1327 205 1331 211
rect 1148 156 1171 161
rect -269 99 -205 102
rect -269 95 -266 99
rect -262 95 -244 99
rect -240 95 -234 99
rect -230 95 -212 99
rect -208 95 -205 99
rect -470 91 -282 94
rect -269 93 -205 95
rect -470 87 -467 91
rect -463 87 -445 91
rect -441 87 -415 91
rect -411 87 -393 91
rect -389 87 -363 91
rect -359 87 -341 91
rect -337 87 -311 91
rect -307 87 -289 91
rect -285 87 -282 91
rect -470 85 -282 87
rect -259 87 -255 93
rect -227 87 -223 93
rect 1148 90 1153 156
rect 1179 152 1183 165
rect 1171 148 1183 152
rect 1201 156 1223 161
rect 1171 143 1175 148
rect 1166 94 1171 99
rect 1179 90 1183 103
rect 1201 90 1206 156
rect 1231 152 1235 165
rect 1283 161 1287 165
rect 1335 161 1339 165
rect 1380 161 1384 173
rect 1412 161 1416 173
rect 1223 148 1235 152
rect 1253 156 1275 161
rect 1283 156 1327 161
rect 1335 156 1372 161
rect 1380 156 1404 161
rect 1412 156 1426 161
rect 1223 143 1227 148
rect 1218 94 1223 99
rect 1231 90 1235 103
rect 1253 90 1258 156
rect 1272 133 1275 138
rect 1283 129 1287 156
rect 1275 98 1279 109
rect 1275 94 1287 98
rect -460 79 -456 85
rect -408 79 -404 85
rect -356 79 -352 85
rect -304 79 -300 85
rect 1148 85 1171 90
rect 1179 85 1223 90
rect 1231 85 1275 90
rect 1179 82 1183 85
rect 1231 82 1235 85
rect 1283 82 1287 94
rect 1305 90 1310 156
rect 1324 133 1327 138
rect 1335 129 1339 156
rect 1380 153 1384 156
rect 1412 153 1416 156
rect 1372 126 1376 133
rect 1404 126 1408 133
rect 1362 124 1426 126
rect 1362 120 1364 124
rect 1368 120 1388 124
rect 1392 120 1396 124
rect 1400 120 1420 124
rect 1424 120 1426 124
rect 1362 118 1426 120
rect 1327 98 1331 109
rect 1327 94 1339 98
rect 1305 85 1327 90
rect 1335 82 1339 94
rect 1171 54 1175 62
rect 1223 54 1227 62
rect 1275 54 1279 62
rect 1327 54 1331 62
rect 1161 53 1349 54
rect 1161 49 1188 53
rect 1192 49 1240 53
rect 1244 49 1292 53
rect 1296 49 1344 53
rect 1348 49 1349 53
rect 1161 48 1349 49
rect -483 30 -460 35
rect -483 -36 -478 30
rect -452 26 -448 39
rect -460 22 -448 26
rect -430 30 -408 35
rect -460 17 -456 22
rect -465 -32 -460 -27
rect -452 -36 -448 -23
rect -430 -36 -425 30
rect -400 26 -396 39
rect -348 35 -344 39
rect -296 35 -292 39
rect -251 35 -247 47
rect -219 35 -215 47
rect 618 39 645 42
rect 618 35 621 39
rect 625 35 638 39
rect 642 35 645 39
rect 1154 35 1161 40
rect 1166 35 1213 40
rect 1218 35 1267 40
rect 1272 35 1319 40
rect -408 22 -396 26
rect -378 30 -356 35
rect -348 30 -304 35
rect -296 30 -259 35
rect -251 30 -227 35
rect -219 30 -205 35
rect 618 33 645 35
rect -408 17 -404 22
rect -413 -32 -408 -27
rect -400 -36 -396 -23
rect -378 -36 -373 30
rect -359 7 -356 12
rect -348 3 -344 30
rect -356 -28 -352 -17
rect -356 -32 -344 -28
rect -483 -41 -460 -36
rect -452 -41 -408 -36
rect -400 -41 -356 -36
rect -452 -44 -448 -41
rect -400 -44 -396 -41
rect -348 -44 -344 -32
rect -326 -36 -321 30
rect -307 7 -304 12
rect -296 3 -292 30
rect -251 27 -247 30
rect -219 27 -215 30
rect -31 26 299 30
rect 304 26 434 30
rect 626 28 630 33
rect 431 20 434 26
rect 515 20 520 22
rect 431 15 520 20
rect 480 11 486 12
rect 480 7 481 11
rect 485 7 486 11
rect -259 0 -255 7
rect -227 0 -223 7
rect 480 4 486 7
rect 515 4 520 15
rect 575 9 584 12
rect 575 5 577 9
rect 581 5 584 9
rect 598 5 611 8
rect 575 4 584 5
rect 480 0 492 4
rect -269 -2 -205 0
rect -269 -6 -267 -2
rect -263 -6 -243 -2
rect -239 -6 -235 -2
rect -231 -6 -211 -2
rect -207 -6 -205 -2
rect -269 -8 -205 -6
rect 480 -10 486 0
rect 570 0 584 4
rect 512 -8 530 -4
rect 575 -8 584 0
rect 480 -14 481 -10
rect 485 -14 486 -10
rect 480 -15 486 -14
rect -304 -28 -300 -17
rect 313 -22 434 -17
rect 515 -18 520 -8
rect 575 -12 577 -8
rect 581 -12 584 -8
rect 575 -15 584 -12
rect 590 -18 594 -15
rect 431 -27 435 -22
rect 544 -22 594 -18
rect 544 -27 548 -22
rect -304 -32 -292 -28
rect 431 -32 548 -27
rect 598 -28 602 -15
rect 605 -22 611 5
rect 634 -22 638 -12
rect 605 -27 626 -22
rect 634 -27 683 -22
rect -326 -41 -304 -36
rect -296 -44 -292 -32
rect 480 -40 486 -39
rect 480 -44 481 -40
rect 485 -44 486 -40
rect 480 -47 486 -44
rect 515 -47 520 -32
rect 575 -42 584 -39
rect 575 -46 577 -42
rect 581 -46 584 -42
rect 575 -47 584 -46
rect 480 -51 492 -47
rect 480 -61 486 -51
rect 570 -51 584 -47
rect 512 -59 530 -55
rect 575 -59 584 -51
rect -460 -72 -456 -64
rect -408 -72 -404 -64
rect -356 -72 -352 -64
rect -304 -72 -300 -64
rect 480 -65 481 -61
rect 485 -65 486 -61
rect 480 -66 486 -65
rect -470 -73 -282 -72
rect -470 -77 -443 -73
rect -439 -77 -391 -73
rect -387 -77 -339 -73
rect -335 -77 -287 -73
rect -283 -77 -282 -73
rect -470 -78 -282 -77
rect 515 -79 520 -59
rect 575 -63 577 -59
rect 581 -63 584 -59
rect 575 -66 584 -63
rect 634 -30 638 -27
rect 590 -79 594 -48
rect 626 -56 630 -50
rect 618 -57 645 -56
rect 618 -61 619 -57
rect 623 -61 640 -57
rect 644 -61 645 -57
rect 618 -62 645 -61
rect 515 -82 594 -79
rect -477 -91 -470 -86
rect -465 -91 -418 -86
rect -413 -91 -364 -86
rect -359 -91 -312 -86
rect 712 -135 739 -132
rect 712 -139 715 -135
rect 719 -139 732 -135
rect 736 -139 739 -135
rect 712 -141 739 -139
rect 720 -146 724 -141
rect 246 -152 273 -149
rect 246 -156 249 -152
rect 253 -156 266 -152
rect 270 -156 273 -152
rect 246 -158 273 -156
rect 254 -163 258 -158
rect 143 -171 148 -169
rect -19 -176 14 -171
rect 19 -176 148 -171
rect 108 -180 114 -179
rect 108 -184 109 -180
rect 113 -184 114 -180
rect 108 -187 114 -184
rect 143 -187 148 -176
rect 203 -182 212 -179
rect 203 -186 205 -182
rect 209 -186 212 -182
rect 226 -186 239 -183
rect 203 -187 212 -186
rect 108 -191 120 -187
rect 108 -201 114 -191
rect 198 -191 212 -187
rect 140 -199 158 -195
rect 203 -199 212 -191
rect 108 -205 109 -201
rect 113 -205 114 -201
rect 108 -206 114 -205
rect 143 -209 148 -199
rect 203 -203 205 -199
rect 209 -203 212 -199
rect 203 -206 212 -203
rect 218 -209 222 -206
rect 172 -213 222 -209
rect 172 -218 176 -213
rect -16 -223 176 -218
rect 226 -219 230 -206
rect 233 -213 239 -186
rect 467 -168 521 -165
rect 467 -172 470 -168
rect 474 -172 487 -168
rect 491 -172 497 -168
rect 501 -172 514 -168
rect 518 -172 521 -168
rect 467 -174 521 -172
rect 262 -213 266 -203
rect 475 -179 479 -174
rect 502 -179 506 -174
rect 233 -218 254 -213
rect 262 -218 308 -213
rect 313 -214 407 -213
rect 313 -218 431 -214
rect -236 -296 -172 -293
rect -236 -300 -233 -296
rect -229 -300 -211 -296
rect -207 -300 -201 -296
rect -197 -300 -179 -296
rect -175 -300 -172 -296
rect -437 -304 -249 -301
rect -236 -302 -172 -300
rect -437 -308 -434 -304
rect -430 -308 -412 -304
rect -408 -308 -382 -304
rect -378 -308 -360 -304
rect -356 -308 -330 -304
rect -326 -308 -308 -304
rect -304 -308 -278 -304
rect -274 -308 -256 -304
rect -252 -308 -249 -304
rect -437 -310 -249 -308
rect -226 -308 -222 -302
rect -194 -308 -190 -302
rect -427 -316 -423 -310
rect -375 -316 -371 -310
rect -323 -316 -319 -310
rect -271 -316 -267 -310
rect -450 -365 -427 -360
rect -450 -431 -445 -365
rect -419 -369 -415 -356
rect -427 -373 -415 -369
rect -397 -365 -375 -360
rect -427 -378 -423 -373
rect -432 -427 -427 -422
rect -419 -431 -415 -418
rect -397 -431 -392 -365
rect -367 -369 -363 -356
rect -315 -360 -311 -356
rect -263 -360 -259 -356
rect -218 -360 -214 -348
rect -186 -360 -182 -348
rect -375 -373 -363 -369
rect -345 -365 -323 -360
rect -315 -365 -271 -360
rect -263 -365 -226 -360
rect -218 -365 -194 -360
rect -186 -365 -172 -360
rect -375 -378 -371 -373
rect -380 -427 -375 -422
rect -367 -431 -363 -418
rect -345 -431 -340 -365
rect -326 -388 -323 -383
rect -315 -392 -311 -365
rect -323 -423 -319 -412
rect -323 -427 -311 -423
rect -450 -436 -427 -431
rect -419 -436 -375 -431
rect -367 -436 -323 -431
rect -419 -439 -415 -436
rect -367 -439 -363 -436
rect -315 -439 -311 -427
rect -293 -431 -288 -365
rect -274 -388 -271 -383
rect -263 -392 -259 -365
rect -218 -368 -214 -365
rect -186 -368 -182 -365
rect -226 -395 -222 -388
rect -194 -395 -190 -388
rect -236 -397 -172 -395
rect -236 -401 -234 -397
rect -230 -401 -210 -397
rect -206 -401 -202 -397
rect -198 -401 -178 -397
rect -174 -401 -172 -397
rect -236 -403 -172 -401
rect -271 -423 -267 -412
rect -271 -427 -259 -423
rect -293 -436 -271 -431
rect -263 -439 -259 -427
rect 69 -438 74 -223
rect 108 -231 114 -230
rect 108 -235 109 -231
rect 113 -235 114 -231
rect 108 -238 114 -235
rect 143 -238 148 -223
rect 203 -233 212 -230
rect 203 -237 205 -233
rect 209 -237 212 -233
rect 203 -238 212 -237
rect 108 -242 120 -238
rect 108 -252 114 -242
rect 198 -242 212 -238
rect 140 -250 158 -246
rect 203 -250 212 -242
rect 108 -256 109 -252
rect 113 -256 114 -252
rect 108 -257 114 -256
rect 143 -270 148 -250
rect 203 -254 205 -250
rect 209 -254 212 -250
rect 203 -257 212 -254
rect 262 -221 266 -218
rect 218 -270 222 -239
rect 254 -247 258 -241
rect 397 -244 431 -218
rect 483 -239 487 -219
rect 510 -239 514 -219
rect 632 -234 720 -229
rect 529 -238 556 -235
rect 483 -243 524 -239
rect 246 -248 273 -247
rect 246 -252 247 -248
rect 251 -252 268 -248
rect 272 -252 273 -248
rect 397 -249 475 -244
rect 397 -250 431 -249
rect 246 -253 273 -252
rect 502 -253 506 -243
rect 143 -273 222 -270
rect 304 -280 407 -279
rect 304 -284 429 -280
rect 163 -296 217 -293
rect 163 -300 166 -296
rect 170 -300 183 -296
rect 187 -300 193 -296
rect 197 -300 210 -296
rect 214 -300 217 -296
rect 163 -302 217 -300
rect 171 -307 175 -302
rect 198 -307 202 -302
rect 399 -310 429 -284
rect 494 -299 498 -293
rect 519 -299 524 -243
rect 529 -242 532 -238
rect 536 -242 549 -238
rect 553 -242 556 -238
rect 529 -244 556 -242
rect 537 -249 541 -244
rect 545 -299 549 -289
rect 574 -299 602 -298
rect 494 -303 508 -299
rect 502 -304 508 -303
rect 519 -304 537 -299
rect 545 -304 602 -299
rect 399 -315 494 -310
rect 502 -318 506 -304
rect 545 -307 549 -304
rect 179 -367 183 -347
rect 206 -367 210 -347
rect 537 -333 541 -327
rect 529 -334 556 -333
rect 529 -338 530 -334
rect 534 -338 551 -334
rect 555 -338 556 -334
rect 529 -339 556 -338
rect 574 -351 602 -304
rect 632 -351 637 -234
rect 728 -238 732 -226
rect 720 -242 732 -238
rect 1640 -238 1704 -235
rect 1640 -242 1643 -238
rect 1647 -242 1665 -238
rect 1669 -242 1675 -238
rect 1679 -242 1697 -238
rect 1701 -242 1704 -238
rect 720 -246 724 -242
rect 1439 -246 1627 -243
rect 1640 -244 1704 -242
rect 1439 -250 1442 -246
rect 1446 -250 1464 -246
rect 1468 -250 1494 -246
rect 1498 -250 1516 -246
rect 1520 -250 1546 -246
rect 1550 -250 1568 -246
rect 1572 -250 1598 -246
rect 1602 -250 1620 -246
rect 1624 -250 1627 -246
rect 1439 -252 1627 -250
rect 1650 -250 1654 -244
rect 1682 -250 1686 -244
rect 1449 -258 1453 -252
rect 1501 -258 1505 -252
rect 1553 -258 1557 -252
rect 1605 -258 1609 -252
rect 761 -272 788 -269
rect 761 -276 764 -272
rect 768 -276 781 -272
rect 785 -276 788 -272
rect 761 -278 788 -276
rect 769 -283 773 -278
rect 574 -356 637 -351
rect 661 -337 705 -332
rect 728 -333 732 -326
rect 777 -333 781 -323
rect 1426 -307 1449 -302
rect 574 -357 602 -356
rect 225 -366 252 -363
rect 494 -364 498 -358
rect 179 -371 220 -367
rect 107 -377 171 -372
rect 198 -381 202 -371
rect 190 -427 194 -421
rect 215 -427 220 -371
rect 225 -370 228 -366
rect 232 -370 245 -366
rect 249 -370 252 -366
rect 486 -365 513 -364
rect 486 -369 487 -365
rect 491 -369 508 -365
rect 512 -369 513 -365
rect 486 -370 513 -369
rect 225 -372 252 -370
rect 233 -377 237 -372
rect 241 -427 245 -417
rect 190 -431 204 -427
rect 198 -432 204 -431
rect 215 -432 233 -427
rect 241 -432 317 -427
rect 322 -428 407 -427
rect 322 -432 432 -428
rect 69 -443 190 -438
rect 198 -446 202 -432
rect 241 -435 245 -432
rect -427 -467 -423 -459
rect -375 -467 -371 -459
rect -323 -467 -319 -459
rect -271 -467 -267 -459
rect -437 -468 -249 -467
rect -437 -472 -410 -468
rect -406 -472 -358 -468
rect -354 -472 -306 -468
rect -302 -472 -254 -468
rect -250 -472 -249 -468
rect -437 -473 -249 -472
rect -444 -486 -437 -481
rect -432 -486 -385 -481
rect -380 -486 -331 -481
rect -326 -486 -279 -481
rect 233 -461 237 -455
rect 403 -456 432 -432
rect 331 -461 391 -456
rect 402 -458 432 -456
rect 402 -459 578 -458
rect 402 -461 637 -459
rect 225 -462 252 -461
rect 225 -466 226 -462
rect 230 -466 247 -462
rect 251 -466 252 -462
rect 225 -467 252 -466
rect 190 -492 194 -486
rect 375 -487 389 -461
rect 403 -463 637 -461
rect 374 -492 556 -487
rect 182 -493 209 -492
rect 182 -497 183 -493
rect 187 -497 204 -493
rect 208 -497 209 -493
rect 374 -495 427 -492
rect 375 -496 389 -495
rect 182 -498 209 -497
rect 525 -539 556 -492
rect 571 -510 637 -463
rect 661 -510 666 -337
rect 728 -338 769 -333
rect 777 -338 865 -333
rect 728 -341 732 -338
rect 777 -341 781 -338
rect 713 -345 750 -341
rect 713 -351 717 -345
rect 746 -351 750 -345
rect 769 -367 773 -361
rect 761 -368 788 -367
rect 705 -377 709 -371
rect 738 -377 742 -371
rect 761 -372 762 -368
rect 766 -372 783 -368
rect 787 -372 788 -368
rect 761 -373 788 -372
rect 697 -378 724 -377
rect 697 -382 698 -378
rect 702 -382 719 -378
rect 723 -382 724 -378
rect 697 -383 724 -382
rect 730 -378 757 -377
rect 730 -382 731 -378
rect 735 -382 752 -378
rect 756 -382 757 -378
rect 730 -383 757 -382
rect 846 -427 865 -338
rect 1114 -348 1141 -345
rect 1114 -352 1117 -348
rect 1121 -352 1134 -348
rect 1138 -352 1141 -348
rect 1114 -354 1141 -352
rect 1122 -359 1126 -354
rect 1011 -367 1016 -365
rect 939 -372 1016 -367
rect 939 -427 944 -372
rect 976 -376 982 -375
rect 976 -380 977 -376
rect 981 -380 982 -376
rect 976 -383 982 -380
rect 1011 -383 1016 -372
rect 1071 -378 1080 -375
rect 1071 -382 1073 -378
rect 1077 -382 1080 -378
rect 1094 -382 1107 -379
rect 1071 -383 1080 -382
rect 976 -387 988 -383
rect 976 -397 982 -387
rect 1066 -387 1080 -383
rect 1008 -395 1026 -391
rect 1071 -395 1080 -387
rect 976 -401 977 -397
rect 981 -401 982 -397
rect 976 -402 982 -401
rect 1011 -405 1016 -395
rect 1071 -399 1073 -395
rect 1077 -399 1080 -395
rect 1071 -402 1080 -399
rect 1086 -405 1090 -402
rect 1040 -409 1090 -405
rect 1040 -414 1044 -409
rect 846 -432 944 -427
rect 953 -419 1044 -414
rect 1094 -415 1098 -402
rect 1101 -409 1107 -382
rect 1426 -373 1431 -307
rect 1457 -311 1461 -298
rect 1449 -315 1461 -311
rect 1479 -307 1501 -302
rect 1449 -320 1453 -315
rect 1444 -369 1449 -364
rect 1457 -373 1461 -360
rect 1479 -373 1484 -307
rect 1509 -311 1513 -298
rect 1561 -302 1565 -298
rect 1613 -302 1617 -298
rect 1658 -302 1662 -290
rect 1690 -302 1694 -290
rect 1501 -315 1513 -311
rect 1531 -307 1553 -302
rect 1561 -307 1605 -302
rect 1613 -307 1650 -302
rect 1658 -307 1682 -302
rect 1690 -307 1704 -302
rect 1501 -320 1505 -315
rect 1496 -369 1501 -364
rect 1509 -373 1513 -360
rect 1531 -373 1536 -307
rect 1550 -330 1553 -325
rect 1561 -334 1565 -307
rect 1553 -365 1557 -354
rect 1553 -369 1565 -365
rect 1426 -378 1449 -373
rect 1457 -378 1501 -373
rect 1509 -378 1553 -373
rect 1457 -381 1461 -378
rect 1509 -381 1513 -378
rect 1561 -381 1565 -369
rect 1583 -373 1588 -307
rect 1602 -330 1605 -325
rect 1613 -334 1617 -307
rect 1658 -310 1662 -307
rect 1690 -310 1694 -307
rect 1650 -337 1654 -330
rect 1682 -337 1686 -330
rect 1640 -339 1704 -337
rect 1640 -343 1642 -339
rect 1646 -343 1666 -339
rect 1670 -343 1674 -339
rect 1678 -343 1698 -339
rect 1702 -343 1704 -339
rect 1640 -345 1704 -343
rect 1605 -365 1609 -354
rect 1605 -369 1617 -365
rect 1583 -378 1605 -373
rect 1613 -381 1617 -369
rect 1130 -409 1134 -399
rect 1449 -409 1453 -401
rect 1501 -409 1505 -401
rect 1553 -409 1557 -401
rect 1605 -409 1609 -401
rect 1101 -414 1122 -409
rect 1130 -414 1172 -409
rect 1439 -410 1627 -409
rect 1439 -414 1466 -410
rect 1470 -414 1518 -410
rect 1522 -414 1570 -410
rect 1574 -414 1622 -410
rect 1626 -414 1627 -410
rect 953 -466 958 -419
rect 976 -427 982 -426
rect 976 -431 977 -427
rect 981 -431 982 -427
rect 976 -434 982 -431
rect 1011 -434 1016 -419
rect 1071 -429 1080 -426
rect 1071 -433 1073 -429
rect 1077 -433 1080 -429
rect 1071 -434 1080 -433
rect 976 -438 988 -434
rect 976 -448 982 -438
rect 1066 -438 1080 -434
rect 1008 -446 1026 -442
rect 1071 -446 1080 -438
rect 976 -452 977 -448
rect 981 -452 982 -448
rect 976 -453 982 -452
rect 842 -484 958 -466
rect 1011 -466 1016 -446
rect 1071 -450 1073 -446
rect 1077 -450 1080 -446
rect 1071 -453 1080 -450
rect 1130 -417 1134 -414
rect 1439 -415 1627 -414
rect 1086 -466 1090 -435
rect 1432 -428 1439 -423
rect 1444 -428 1491 -423
rect 1496 -428 1545 -423
rect 1550 -428 1597 -423
rect 1122 -443 1126 -437
rect 1114 -444 1141 -443
rect 1114 -448 1115 -444
rect 1119 -448 1136 -444
rect 1140 -448 1141 -444
rect 1114 -449 1141 -448
rect 1011 -469 1090 -466
rect 571 -515 666 -510
rect 841 -488 958 -484
rect 841 -539 864 -488
rect 953 -489 958 -488
rect 525 -544 865 -539
rect 525 -545 583 -544
rect 841 -545 864 -544
rect 1193 -616 1220 -613
rect 1193 -620 1196 -616
rect 1200 -620 1213 -616
rect 1217 -620 1220 -616
rect 967 -624 994 -621
rect 1193 -622 1220 -620
rect 967 -628 970 -624
rect 974 -628 987 -624
rect 991 -628 994 -624
rect 298 -635 303 -634
rect 925 -635 930 -629
rect 967 -630 994 -628
rect 1201 -627 1205 -622
rect 298 -646 930 -635
rect -345 -675 -281 -672
rect -345 -679 -342 -675
rect -338 -679 -320 -675
rect -316 -679 -310 -675
rect -306 -679 -288 -675
rect -284 -679 -281 -675
rect -546 -683 -358 -680
rect -345 -681 -281 -679
rect -546 -687 -543 -683
rect -539 -687 -521 -683
rect -517 -687 -491 -683
rect -487 -687 -469 -683
rect -465 -687 -439 -683
rect -435 -687 -417 -683
rect -413 -687 -387 -683
rect -383 -687 -365 -683
rect -361 -687 -358 -683
rect -546 -689 -358 -687
rect -335 -687 -331 -681
rect -303 -687 -299 -681
rect -536 -695 -532 -689
rect -484 -695 -480 -689
rect -432 -695 -428 -689
rect -380 -695 -376 -689
rect 298 -709 303 -646
rect 568 -657 622 -654
rect 568 -661 571 -657
rect 575 -661 588 -657
rect 592 -661 598 -657
rect 602 -661 615 -657
rect 619 -661 622 -657
rect 568 -663 622 -661
rect 576 -668 580 -663
rect 603 -668 607 -663
rect 298 -717 303 -714
rect -559 -744 -536 -739
rect -559 -810 -554 -744
rect -528 -748 -524 -735
rect -536 -752 -524 -748
rect -506 -744 -484 -739
rect -536 -757 -532 -752
rect -541 -806 -536 -801
rect -528 -810 -524 -797
rect -506 -810 -501 -744
rect -476 -748 -472 -735
rect -424 -739 -420 -735
rect -372 -739 -368 -735
rect -327 -739 -323 -727
rect -295 -739 -291 -727
rect 584 -728 588 -708
rect 611 -728 615 -708
rect 925 -718 930 -646
rect 975 -635 979 -630
rect 925 -723 975 -718
rect 630 -727 657 -724
rect 983 -727 987 -715
rect 584 -732 625 -728
rect 285 -738 576 -733
rect -484 -752 -472 -748
rect -454 -744 -432 -739
rect -424 -744 -380 -739
rect -372 -744 -335 -739
rect -327 -744 -303 -739
rect -295 -744 -281 -739
rect 603 -742 607 -732
rect -484 -757 -480 -752
rect -489 -806 -484 -801
rect -476 -810 -472 -797
rect -454 -810 -449 -744
rect -435 -767 -432 -762
rect -424 -771 -420 -744
rect -432 -802 -428 -791
rect -432 -806 -420 -802
rect -559 -815 -536 -810
rect -528 -815 -484 -810
rect -476 -815 -432 -810
rect -528 -818 -524 -815
rect -476 -818 -472 -815
rect -424 -818 -420 -806
rect -402 -810 -397 -744
rect -383 -767 -380 -762
rect -372 -771 -368 -744
rect -327 -747 -323 -744
rect -295 -747 -291 -744
rect -335 -774 -331 -767
rect -303 -774 -299 -767
rect -345 -776 -281 -774
rect -345 -780 -343 -776
rect -339 -780 -319 -776
rect -315 -780 -311 -776
rect -307 -780 -287 -776
rect -283 -780 -281 -776
rect -345 -782 -281 -780
rect 197 -788 224 -785
rect -380 -802 -376 -791
rect 197 -792 200 -788
rect 204 -792 217 -788
rect 221 -792 224 -788
rect 595 -788 599 -782
rect 620 -788 625 -732
rect 630 -731 633 -727
rect 637 -731 650 -727
rect 654 -731 657 -727
rect 630 -733 657 -731
rect 975 -731 987 -727
rect 1085 -711 1122 -707
rect 1167 -711 1201 -710
rect 1085 -715 1201 -711
rect 1085 -724 1174 -715
rect 1209 -719 1213 -707
rect 1201 -723 1213 -719
rect 638 -738 642 -733
rect 975 -735 979 -731
rect 646 -788 650 -778
rect 595 -792 609 -788
rect 197 -794 224 -792
rect 603 -793 609 -792
rect 620 -793 638 -788
rect 646 -793 953 -788
rect 205 -799 209 -794
rect -380 -806 -368 -802
rect -402 -815 -380 -810
rect -372 -818 -368 -806
rect 94 -807 99 -805
rect -68 -812 -35 -807
rect -30 -812 99 -807
rect 59 -816 65 -815
rect 59 -820 60 -816
rect 64 -820 65 -816
rect 59 -823 65 -820
rect 94 -823 99 -812
rect 154 -818 163 -815
rect 154 -822 156 -818
rect 160 -822 163 -818
rect 177 -822 190 -819
rect 154 -823 163 -822
rect 59 -827 71 -823
rect 59 -837 65 -827
rect 149 -827 163 -823
rect 91 -835 109 -831
rect 154 -835 163 -827
rect -536 -846 -532 -838
rect -484 -846 -480 -838
rect -432 -846 -428 -838
rect -380 -846 -376 -838
rect 59 -841 60 -837
rect 64 -841 65 -837
rect 59 -842 65 -841
rect 94 -845 99 -835
rect 154 -839 156 -835
rect 160 -839 163 -835
rect 154 -842 163 -839
rect 169 -845 173 -842
rect -546 -847 -358 -846
rect -546 -851 -519 -847
rect -515 -851 -467 -847
rect -463 -851 -415 -847
rect -411 -851 -363 -847
rect -359 -851 -358 -847
rect 123 -849 173 -845
rect -546 -852 -358 -851
rect 123 -854 127 -849
rect -65 -859 127 -854
rect 177 -855 181 -842
rect 184 -849 190 -822
rect 213 -849 217 -839
rect 530 -804 595 -799
rect 530 -849 535 -804
rect 603 -807 607 -793
rect 646 -796 650 -793
rect 184 -854 205 -849
rect 213 -854 289 -849
rect 294 -854 535 -849
rect 638 -822 642 -816
rect 948 -821 953 -793
rect 1016 -761 1043 -758
rect 1016 -765 1019 -761
rect 1023 -765 1036 -761
rect 1040 -765 1043 -761
rect 1016 -767 1043 -765
rect 1024 -772 1028 -767
rect 630 -823 657 -822
rect 630 -827 631 -823
rect 635 -827 652 -823
rect 656 -827 657 -823
rect 948 -826 960 -821
rect 983 -822 987 -815
rect 1032 -822 1036 -812
rect 1085 -821 1122 -724
rect 1201 -727 1205 -723
rect 1242 -753 1269 -750
rect 1242 -757 1245 -753
rect 1249 -757 1262 -753
rect 1266 -757 1269 -753
rect 1242 -759 1269 -757
rect 1250 -764 1254 -759
rect 1468 -793 1495 -790
rect 1468 -797 1471 -793
rect 1475 -797 1488 -793
rect 1492 -797 1495 -793
rect 1468 -799 1495 -797
rect 1951 -793 2015 -790
rect 1951 -797 1954 -793
rect 1958 -797 1976 -793
rect 1980 -797 1986 -793
rect 1990 -797 2008 -793
rect 2012 -797 2015 -793
rect 1061 -822 1122 -821
rect 630 -828 657 -827
rect 983 -827 1024 -822
rect 1032 -827 1122 -822
rect 983 -830 987 -827
rect 1032 -830 1036 -827
rect 1061 -828 1122 -827
rect 1149 -818 1186 -813
rect 1209 -814 1213 -807
rect 1258 -814 1262 -804
rect 1476 -804 1480 -799
rect 1750 -801 1938 -798
rect 1951 -799 2015 -797
rect 1365 -812 1370 -810
rect 1311 -814 1370 -812
rect 968 -834 1005 -830
rect 968 -840 972 -834
rect 1001 -840 1005 -834
rect 595 -853 599 -847
rect 587 -854 614 -853
rect -553 -865 -546 -860
rect -541 -865 -494 -860
rect -489 -865 -440 -860
rect -435 -865 -388 -860
rect -269 -1028 -205 -1025
rect -269 -1032 -266 -1028
rect -262 -1032 -244 -1028
rect -240 -1032 -234 -1028
rect -230 -1032 -212 -1028
rect -208 -1032 -205 -1028
rect -470 -1036 -282 -1033
rect -269 -1034 -205 -1032
rect -470 -1040 -467 -1036
rect -463 -1040 -445 -1036
rect -441 -1040 -415 -1036
rect -411 -1040 -393 -1036
rect -389 -1040 -363 -1036
rect -359 -1040 -341 -1036
rect -337 -1040 -311 -1036
rect -307 -1040 -289 -1036
rect -285 -1040 -282 -1036
rect -470 -1042 -282 -1040
rect -259 -1040 -255 -1034
rect -227 -1040 -223 -1034
rect -460 -1048 -456 -1042
rect -408 -1048 -404 -1042
rect -356 -1048 -352 -1042
rect -304 -1048 -300 -1042
rect 20 -1074 25 -859
rect 59 -867 65 -866
rect 59 -871 60 -867
rect 64 -871 65 -867
rect 59 -874 65 -871
rect 94 -874 99 -859
rect 154 -869 163 -866
rect 154 -873 156 -869
rect 160 -873 163 -869
rect 154 -874 163 -873
rect 59 -878 71 -874
rect 59 -888 65 -878
rect 149 -878 163 -874
rect 91 -886 109 -882
rect 154 -886 163 -878
rect 59 -892 60 -888
rect 64 -892 65 -888
rect 59 -893 65 -892
rect 94 -906 99 -886
rect 154 -890 156 -886
rect 160 -890 163 -886
rect 154 -893 163 -890
rect 213 -857 217 -854
rect 169 -906 173 -875
rect 587 -858 588 -854
rect 592 -858 609 -854
rect 613 -858 614 -854
rect 587 -859 614 -858
rect 1024 -856 1028 -850
rect 1016 -857 1043 -856
rect 960 -866 964 -860
rect 993 -866 997 -860
rect 1016 -861 1017 -857
rect 1021 -861 1038 -857
rect 1042 -861 1043 -857
rect 1016 -862 1043 -861
rect 952 -867 979 -866
rect 952 -871 953 -867
rect 957 -871 974 -867
rect 978 -871 979 -867
rect 952 -872 979 -871
rect 985 -867 1012 -866
rect 985 -871 986 -867
rect 990 -871 1007 -867
rect 1011 -871 1012 -867
rect 985 -872 1012 -871
rect 205 -883 209 -877
rect 197 -884 224 -883
rect 197 -888 198 -884
rect 202 -888 219 -884
rect 223 -888 224 -884
rect 197 -889 224 -888
rect 94 -909 173 -906
rect 491 -902 545 -899
rect 491 -906 494 -902
rect 498 -906 511 -902
rect 515 -906 521 -902
rect 525 -906 538 -902
rect 542 -906 545 -902
rect 491 -908 545 -906
rect 709 -902 763 -899
rect 709 -906 712 -902
rect 716 -906 729 -902
rect 733 -906 739 -902
rect 743 -906 756 -902
rect 760 -906 763 -902
rect 709 -908 763 -906
rect 499 -913 503 -908
rect 526 -913 530 -908
rect 717 -913 721 -908
rect 744 -913 748 -908
rect 114 -932 168 -929
rect 114 -936 117 -932
rect 121 -936 134 -932
rect 138 -936 144 -932
rect 148 -936 161 -932
rect 165 -936 168 -932
rect 114 -938 168 -936
rect 122 -943 126 -938
rect 149 -943 153 -938
rect 507 -973 511 -953
rect 534 -973 538 -953
rect 553 -972 580 -969
rect 507 -977 548 -973
rect 267 -983 499 -978
rect 130 -1003 134 -983
rect 157 -1003 161 -983
rect 526 -987 530 -977
rect 276 -995 487 -990
rect 176 -1002 203 -999
rect 130 -1007 171 -1003
rect 58 -1013 122 -1008
rect 149 -1017 153 -1007
rect 141 -1063 145 -1057
rect 166 -1063 171 -1007
rect 176 -1006 179 -1002
rect 183 -1006 196 -1002
rect 200 -1006 203 -1002
rect 176 -1008 203 -1006
rect 184 -1013 188 -1008
rect 482 -1044 487 -995
rect 518 -1033 522 -1027
rect 543 -1033 548 -977
rect 553 -976 556 -972
rect 560 -976 573 -972
rect 577 -976 580 -972
rect 553 -978 580 -976
rect 725 -973 729 -953
rect 752 -973 756 -953
rect 771 -972 798 -969
rect 725 -977 766 -973
rect 673 -978 705 -977
rect 561 -983 565 -978
rect 613 -983 717 -978
rect 569 -1033 573 -1023
rect 613 -1033 618 -983
rect 744 -987 748 -977
rect 518 -1037 532 -1033
rect 526 -1038 532 -1037
rect 543 -1038 561 -1033
rect 569 -1038 618 -1033
rect 736 -1033 740 -1027
rect 761 -1033 766 -977
rect 771 -976 774 -972
rect 778 -976 791 -972
rect 795 -976 798 -972
rect 771 -978 798 -976
rect 779 -983 783 -978
rect 787 -1033 791 -1023
rect 1149 -1032 1168 -818
rect 1209 -819 1250 -814
rect 1258 -817 1370 -814
rect 1258 -819 1316 -817
rect 1209 -822 1213 -819
rect 1258 -822 1262 -819
rect 1311 -820 1316 -819
rect 1194 -826 1231 -822
rect 1194 -832 1198 -826
rect 1227 -832 1231 -826
rect 1330 -821 1336 -820
rect 1330 -825 1331 -821
rect 1335 -825 1336 -821
rect 1330 -828 1336 -825
rect 1365 -828 1370 -817
rect 1425 -823 1434 -820
rect 1425 -827 1427 -823
rect 1431 -827 1434 -823
rect 1448 -827 1461 -824
rect 1425 -828 1434 -827
rect 1330 -832 1342 -828
rect 1330 -842 1336 -832
rect 1420 -832 1434 -828
rect 1362 -840 1380 -836
rect 1425 -840 1434 -832
rect 1250 -848 1254 -842
rect 1330 -846 1331 -842
rect 1335 -846 1336 -842
rect 1330 -847 1336 -846
rect 1242 -849 1269 -848
rect 1186 -858 1190 -852
rect 1219 -858 1223 -852
rect 1242 -853 1243 -849
rect 1247 -853 1264 -849
rect 1268 -853 1269 -849
rect 1242 -854 1269 -853
rect 1365 -850 1370 -840
rect 1425 -844 1427 -840
rect 1431 -844 1434 -840
rect 1425 -847 1434 -844
rect 1440 -850 1444 -847
rect 1394 -854 1444 -850
rect 1178 -859 1205 -858
rect 1178 -863 1179 -859
rect 1183 -863 1200 -859
rect 1204 -863 1205 -859
rect 1178 -864 1205 -863
rect 1211 -859 1238 -858
rect 1394 -859 1398 -854
rect 1211 -863 1212 -859
rect 1216 -863 1233 -859
rect 1237 -863 1238 -859
rect 1211 -864 1238 -863
rect 1307 -864 1398 -859
rect 1448 -860 1452 -847
rect 1455 -854 1461 -827
rect 1750 -805 1753 -801
rect 1757 -805 1775 -801
rect 1779 -805 1805 -801
rect 1809 -805 1827 -801
rect 1831 -805 1857 -801
rect 1861 -805 1879 -801
rect 1883 -805 1909 -801
rect 1913 -805 1931 -801
rect 1935 -805 1938 -801
rect 1750 -807 1938 -805
rect 1961 -805 1965 -799
rect 1993 -805 1997 -799
rect 1484 -854 1488 -844
rect 1760 -813 1764 -807
rect 1812 -813 1816 -807
rect 1864 -813 1868 -807
rect 1916 -813 1920 -807
rect 1455 -859 1476 -854
rect 1484 -859 1495 -854
rect 1060 -1033 1168 -1032
rect 736 -1037 750 -1033
rect 744 -1038 750 -1037
rect 761 -1038 779 -1033
rect 787 -1038 1168 -1033
rect 482 -1049 518 -1044
rect 526 -1052 530 -1038
rect 569 -1041 573 -1038
rect 192 -1063 196 -1053
rect 141 -1067 155 -1063
rect 149 -1068 155 -1067
rect 166 -1068 184 -1063
rect 192 -1068 298 -1063
rect 303 -1068 327 -1063
rect 20 -1079 141 -1074
rect -483 -1097 -460 -1092
rect -483 -1163 -478 -1097
rect -452 -1101 -448 -1088
rect -460 -1105 -448 -1101
rect -430 -1097 -408 -1092
rect -460 -1110 -456 -1105
rect -465 -1159 -460 -1154
rect -452 -1163 -448 -1150
rect -430 -1163 -425 -1097
rect -400 -1101 -396 -1088
rect -348 -1092 -344 -1088
rect -296 -1092 -292 -1088
rect -251 -1092 -247 -1080
rect -219 -1092 -215 -1080
rect 149 -1082 153 -1068
rect 192 -1071 196 -1068
rect -408 -1105 -396 -1101
rect -378 -1097 -356 -1092
rect -348 -1097 -304 -1092
rect -296 -1097 -259 -1092
rect -251 -1097 -227 -1092
rect -219 -1097 -205 -1092
rect -408 -1110 -404 -1105
rect -413 -1159 -408 -1154
rect -400 -1163 -396 -1150
rect -378 -1163 -373 -1097
rect -359 -1120 -356 -1115
rect -348 -1124 -344 -1097
rect -356 -1155 -352 -1144
rect -356 -1159 -344 -1155
rect -483 -1168 -460 -1163
rect -452 -1168 -408 -1163
rect -400 -1168 -356 -1163
rect -452 -1171 -448 -1168
rect -400 -1171 -396 -1168
rect -348 -1171 -344 -1159
rect -326 -1163 -321 -1097
rect -307 -1120 -304 -1115
rect -296 -1124 -292 -1097
rect -251 -1100 -247 -1097
rect -219 -1100 -215 -1097
rect -259 -1127 -255 -1120
rect -227 -1127 -223 -1120
rect 184 -1097 188 -1091
rect 629 -1049 736 -1044
rect 561 -1067 565 -1061
rect 553 -1068 580 -1067
rect 553 -1072 554 -1068
rect 558 -1072 575 -1068
rect 579 -1072 580 -1068
rect 553 -1073 580 -1072
rect 176 -1098 203 -1097
rect 518 -1098 522 -1092
rect 176 -1102 177 -1098
rect 181 -1102 198 -1098
rect 202 -1102 203 -1098
rect 176 -1103 203 -1102
rect 510 -1099 537 -1098
rect 510 -1103 511 -1099
rect 515 -1103 532 -1099
rect 536 -1103 537 -1099
rect 510 -1104 537 -1103
rect 629 -1116 634 -1049
rect 744 -1052 748 -1038
rect 787 -1041 791 -1038
rect 1060 -1039 1168 -1038
rect 1235 -887 1241 -886
rect 1307 -887 1318 -864
rect 1235 -892 1318 -887
rect 779 -1067 783 -1061
rect 771 -1068 798 -1067
rect 771 -1072 772 -1068
rect 776 -1072 793 -1068
rect 797 -1072 798 -1068
rect 771 -1073 798 -1072
rect 736 -1098 740 -1092
rect 728 -1099 755 -1098
rect 728 -1103 729 -1099
rect 733 -1103 750 -1099
rect 754 -1103 755 -1099
rect 728 -1104 755 -1103
rect 294 -1121 634 -1116
rect -269 -1129 -205 -1127
rect 141 -1128 145 -1122
rect 1061 -1128 1177 -1127
rect 1235 -1128 1241 -892
rect 1307 -893 1318 -892
rect 1330 -872 1336 -871
rect 1330 -876 1331 -872
rect 1335 -876 1336 -872
rect 1330 -879 1336 -876
rect 1365 -879 1370 -864
rect 1425 -874 1434 -871
rect 1425 -878 1427 -874
rect 1431 -878 1434 -874
rect 1425 -879 1434 -878
rect 1330 -883 1342 -879
rect 1330 -893 1336 -883
rect 1420 -883 1434 -879
rect 1362 -891 1380 -887
rect 1425 -891 1434 -883
rect 1330 -897 1331 -893
rect 1335 -897 1336 -893
rect 1330 -898 1336 -897
rect 1365 -911 1370 -891
rect 1425 -895 1427 -891
rect 1431 -895 1434 -891
rect 1425 -898 1434 -895
rect 1484 -862 1488 -859
rect 1440 -911 1444 -880
rect 1737 -862 1760 -857
rect 1476 -888 1480 -882
rect 1468 -889 1495 -888
rect 1468 -893 1469 -889
rect 1473 -893 1490 -889
rect 1494 -893 1495 -889
rect 1468 -894 1495 -893
rect 1365 -914 1444 -911
rect 1737 -928 1742 -862
rect 1768 -866 1772 -853
rect 1760 -870 1772 -866
rect 1790 -862 1812 -857
rect 1760 -875 1764 -870
rect 1755 -924 1760 -919
rect 1768 -928 1772 -915
rect 1790 -928 1795 -862
rect 1820 -866 1824 -853
rect 1872 -857 1876 -853
rect 1924 -857 1928 -853
rect 1969 -857 1973 -845
rect 2001 -857 2005 -845
rect 1812 -870 1824 -866
rect 1842 -862 1864 -857
rect 1872 -862 1916 -857
rect 1924 -862 1961 -857
rect 1969 -862 1993 -857
rect 2001 -862 2015 -857
rect 1812 -875 1816 -870
rect 1807 -924 1812 -919
rect 1820 -928 1824 -915
rect 1842 -928 1847 -862
rect 1861 -885 1864 -880
rect 1872 -889 1876 -862
rect 1864 -920 1868 -909
rect 1864 -924 1876 -920
rect 1737 -933 1760 -928
rect 1768 -933 1812 -928
rect 1820 -933 1864 -928
rect 1768 -936 1772 -933
rect 1820 -936 1824 -933
rect 1872 -936 1876 -924
rect 1894 -928 1899 -862
rect 1913 -885 1916 -880
rect 1924 -889 1928 -862
rect 1969 -865 1973 -862
rect 2001 -865 2005 -862
rect 1961 -892 1965 -885
rect 1993 -892 1997 -885
rect 1951 -894 2015 -892
rect 1951 -898 1953 -894
rect 1957 -898 1977 -894
rect 1981 -898 1985 -894
rect 1989 -898 2009 -894
rect 2013 -898 2015 -894
rect 1951 -900 2015 -898
rect 1916 -920 1920 -909
rect 1916 -924 1928 -920
rect 1894 -933 1916 -928
rect 1924 -936 1928 -924
rect 1760 -964 1764 -956
rect 1812 -964 1816 -956
rect 1864 -964 1868 -956
rect 1916 -964 1920 -956
rect 1750 -965 1938 -964
rect 1750 -969 1777 -965
rect 1781 -969 1829 -965
rect 1833 -969 1881 -965
rect 1885 -969 1933 -965
rect 1937 -969 1938 -965
rect 1750 -970 1938 -969
rect 1743 -983 1750 -978
rect 1755 -983 1802 -978
rect 1807 -983 1856 -978
rect 1861 -983 1908 -978
rect -269 -1133 -267 -1129
rect -263 -1133 -243 -1129
rect -239 -1133 -235 -1129
rect -231 -1133 -211 -1129
rect -207 -1133 -205 -1129
rect -269 -1135 -205 -1133
rect 133 -1129 160 -1128
rect 133 -1133 134 -1129
rect 138 -1133 155 -1129
rect 159 -1133 160 -1129
rect 133 -1134 160 -1133
rect 1061 -1134 1241 -1128
rect 1061 -1138 1177 -1134
rect 307 -1144 1177 -1138
rect -304 -1155 -300 -1144
rect 307 -1149 313 -1144
rect 1061 -1145 1177 -1144
rect 312 -1155 313 -1149
rect -304 -1159 -292 -1155
rect -326 -1168 -304 -1163
rect -296 -1171 -292 -1159
rect 307 -1163 313 -1155
rect 316 -1157 390 -1155
rect 316 -1160 507 -1157
rect 316 -1164 321 -1160
rect 316 -1172 321 -1169
rect 382 -1181 507 -1160
rect 382 -1186 1012 -1181
rect -460 -1199 -456 -1191
rect -408 -1199 -404 -1191
rect -356 -1199 -352 -1191
rect -304 -1199 -300 -1191
rect -470 -1200 -282 -1199
rect -470 -1204 -443 -1200
rect -439 -1204 -391 -1200
rect -387 -1204 -339 -1200
rect -335 -1204 -287 -1200
rect -283 -1204 -282 -1200
rect -470 -1205 -282 -1204
rect -477 -1218 -470 -1213
rect -465 -1218 -418 -1213
rect -413 -1218 -364 -1213
rect -359 -1218 -312 -1213
rect 566 -1220 620 -1217
rect 566 -1224 569 -1220
rect 573 -1224 586 -1220
rect 590 -1224 596 -1220
rect 600 -1224 613 -1220
rect 617 -1224 620 -1220
rect 566 -1226 620 -1224
rect 574 -1231 578 -1226
rect 601 -1231 605 -1226
rect 312 -1275 504 -1270
rect 386 -1296 504 -1275
rect 582 -1291 586 -1271
rect 609 -1291 613 -1271
rect 1007 -1261 1012 -1186
rect 1007 -1263 1081 -1261
rect 1007 -1272 1088 -1263
rect 628 -1290 655 -1287
rect 582 -1295 623 -1291
rect 386 -1301 574 -1296
rect 386 -1302 504 -1301
rect 601 -1305 605 -1295
rect 303 -1338 390 -1336
rect 303 -1341 508 -1338
rect -278 -1356 -214 -1353
rect -278 -1360 -275 -1356
rect -271 -1360 -253 -1356
rect -249 -1360 -243 -1356
rect -239 -1360 -221 -1356
rect -217 -1360 -214 -1356
rect -479 -1364 -291 -1361
rect -278 -1362 -214 -1360
rect 385 -1362 508 -1341
rect 593 -1351 597 -1345
rect 618 -1351 623 -1295
rect 628 -1294 631 -1290
rect 635 -1294 648 -1290
rect 652 -1294 655 -1290
rect 628 -1296 655 -1294
rect 636 -1301 640 -1296
rect 644 -1351 648 -1341
rect 593 -1355 607 -1351
rect 601 -1356 607 -1355
rect 618 -1356 636 -1351
rect 644 -1352 657 -1351
rect 644 -1353 951 -1352
rect 644 -1356 988 -1353
rect -479 -1368 -476 -1364
rect -472 -1368 -454 -1364
rect -450 -1368 -424 -1364
rect -420 -1368 -402 -1364
rect -398 -1368 -372 -1364
rect -368 -1368 -350 -1364
rect -346 -1368 -320 -1364
rect -316 -1368 -298 -1364
rect -294 -1368 -291 -1364
rect -479 -1370 -291 -1368
rect -268 -1368 -264 -1362
rect -236 -1368 -232 -1362
rect 385 -1366 593 -1362
rect 499 -1367 593 -1366
rect -469 -1376 -465 -1370
rect -417 -1376 -413 -1370
rect -365 -1376 -361 -1370
rect -313 -1376 -309 -1370
rect 601 -1370 605 -1356
rect 644 -1359 648 -1356
rect 651 -1357 988 -1356
rect -492 -1425 -469 -1420
rect -492 -1491 -487 -1425
rect -461 -1429 -457 -1416
rect -469 -1433 -457 -1429
rect -439 -1425 -417 -1420
rect -469 -1438 -465 -1433
rect -474 -1487 -469 -1482
rect -461 -1491 -457 -1478
rect -439 -1491 -434 -1425
rect -409 -1429 -405 -1416
rect -357 -1420 -353 -1416
rect -305 -1420 -301 -1416
rect -260 -1420 -256 -1408
rect -228 -1420 -224 -1408
rect 636 -1385 640 -1379
rect 628 -1386 655 -1385
rect 628 -1390 629 -1386
rect 633 -1390 650 -1386
rect 654 -1390 655 -1386
rect 628 -1391 655 -1390
rect 593 -1416 597 -1410
rect 585 -1417 612 -1416
rect -417 -1433 -405 -1429
rect -387 -1425 -365 -1420
rect -357 -1425 -313 -1420
rect -305 -1425 -268 -1420
rect -260 -1425 -236 -1420
rect -228 -1425 -214 -1420
rect 585 -1421 586 -1417
rect 590 -1421 607 -1417
rect 611 -1421 612 -1417
rect 585 -1422 612 -1421
rect -417 -1438 -413 -1433
rect -422 -1487 -417 -1482
rect -409 -1491 -405 -1478
rect -387 -1491 -382 -1425
rect -368 -1448 -365 -1443
rect -357 -1452 -353 -1425
rect -365 -1483 -361 -1472
rect -365 -1487 -353 -1483
rect -492 -1496 -469 -1491
rect -461 -1496 -417 -1491
rect -409 -1496 -365 -1491
rect -461 -1499 -457 -1496
rect -409 -1499 -405 -1496
rect -357 -1499 -353 -1487
rect -335 -1491 -330 -1425
rect -316 -1448 -313 -1443
rect -305 -1452 -301 -1425
rect -260 -1428 -256 -1425
rect -228 -1428 -224 -1425
rect 206 -1448 233 -1445
rect -268 -1455 -264 -1448
rect -236 -1455 -232 -1448
rect 206 -1452 209 -1448
rect 213 -1452 226 -1448
rect 230 -1452 233 -1448
rect 206 -1454 233 -1452
rect 803 -1450 857 -1447
rect 803 -1454 806 -1450
rect 810 -1454 823 -1450
rect 827 -1454 833 -1450
rect 837 -1454 850 -1450
rect 854 -1454 857 -1450
rect -278 -1457 -214 -1455
rect -278 -1461 -276 -1457
rect -272 -1461 -252 -1457
rect -248 -1461 -244 -1457
rect -240 -1461 -220 -1457
rect -216 -1461 -214 -1457
rect 214 -1459 218 -1454
rect 803 -1456 857 -1454
rect -278 -1463 -214 -1461
rect 103 -1467 108 -1465
rect -59 -1472 -26 -1467
rect -21 -1472 108 -1467
rect -313 -1483 -309 -1472
rect 68 -1476 74 -1475
rect 68 -1480 69 -1476
rect 73 -1480 74 -1476
rect 68 -1483 74 -1480
rect 103 -1483 108 -1472
rect 163 -1478 172 -1475
rect 163 -1482 165 -1478
rect 169 -1482 172 -1478
rect 186 -1482 199 -1479
rect 163 -1483 172 -1482
rect -313 -1487 -301 -1483
rect -335 -1496 -313 -1491
rect -305 -1499 -301 -1487
rect 68 -1487 80 -1483
rect 68 -1497 74 -1487
rect 158 -1487 172 -1483
rect 100 -1495 118 -1491
rect 163 -1495 172 -1487
rect 68 -1501 69 -1497
rect 73 -1501 74 -1497
rect 68 -1502 74 -1501
rect 103 -1505 108 -1495
rect 163 -1499 165 -1495
rect 169 -1499 172 -1495
rect 163 -1502 172 -1499
rect 178 -1505 182 -1502
rect 132 -1509 182 -1505
rect 132 -1514 136 -1509
rect -56 -1519 136 -1514
rect 186 -1515 190 -1502
rect 193 -1509 199 -1482
rect 222 -1509 226 -1499
rect 811 -1461 815 -1456
rect 838 -1461 842 -1456
rect 567 -1503 621 -1500
rect 567 -1507 570 -1503
rect 574 -1507 587 -1503
rect 591 -1507 597 -1503
rect 601 -1507 614 -1503
rect 618 -1507 621 -1503
rect 567 -1509 621 -1507
rect 193 -1514 214 -1509
rect 222 -1514 307 -1509
rect 312 -1514 341 -1509
rect 575 -1514 579 -1509
rect 602 -1514 606 -1509
rect -469 -1527 -465 -1519
rect -417 -1527 -413 -1519
rect -365 -1527 -361 -1519
rect -313 -1527 -309 -1519
rect -479 -1528 -291 -1527
rect -479 -1532 -452 -1528
rect -448 -1532 -400 -1528
rect -396 -1532 -348 -1528
rect -344 -1532 -296 -1528
rect -292 -1532 -291 -1528
rect -479 -1533 -291 -1532
rect -486 -1546 -479 -1541
rect -474 -1546 -427 -1541
rect -422 -1546 -373 -1541
rect -368 -1546 -321 -1541
rect -294 -1734 -230 -1731
rect -294 -1738 -291 -1734
rect -287 -1738 -269 -1734
rect -265 -1738 -259 -1734
rect -255 -1738 -237 -1734
rect -233 -1738 -230 -1734
rect -495 -1742 -307 -1739
rect -294 -1740 -230 -1738
rect 29 -1734 34 -1519
rect 68 -1527 74 -1526
rect 68 -1531 69 -1527
rect 73 -1531 74 -1527
rect 68 -1534 74 -1531
rect 103 -1534 108 -1519
rect 163 -1529 172 -1526
rect 163 -1533 165 -1529
rect 169 -1533 172 -1529
rect 163 -1534 172 -1533
rect 68 -1538 80 -1534
rect 68 -1548 74 -1538
rect 158 -1538 172 -1534
rect 100 -1546 118 -1542
rect 163 -1546 172 -1538
rect 68 -1552 69 -1548
rect 73 -1552 74 -1548
rect 68 -1553 74 -1552
rect 103 -1566 108 -1546
rect 163 -1550 165 -1546
rect 169 -1550 172 -1546
rect 163 -1553 172 -1550
rect 222 -1517 226 -1514
rect 178 -1566 182 -1535
rect 214 -1543 218 -1537
rect 206 -1544 233 -1543
rect 206 -1548 207 -1544
rect 211 -1548 228 -1544
rect 232 -1548 233 -1544
rect 206 -1549 233 -1548
rect 312 -1554 390 -1553
rect 819 -1521 823 -1501
rect 846 -1521 850 -1501
rect 940 -1495 988 -1357
rect 1066 -1391 1088 -1272
rect 1146 -1297 1173 -1294
rect 1146 -1301 1149 -1297
rect 1153 -1301 1166 -1297
rect 1170 -1301 1173 -1297
rect 1146 -1303 1173 -1301
rect 1154 -1308 1158 -1303
rect 1063 -1396 1154 -1391
rect 1162 -1400 1166 -1388
rect 1154 -1404 1166 -1400
rect 1154 -1408 1158 -1404
rect 1195 -1434 1222 -1431
rect 1195 -1438 1198 -1434
rect 1202 -1438 1215 -1434
rect 1219 -1438 1222 -1434
rect 1195 -1440 1222 -1438
rect 1203 -1445 1207 -1440
rect 1306 -1461 1333 -1458
rect 1306 -1465 1309 -1461
rect 1313 -1465 1326 -1461
rect 1330 -1465 1333 -1461
rect 1306 -1467 1333 -1465
rect 1063 -1495 1139 -1494
rect 940 -1499 1139 -1495
rect 1162 -1495 1166 -1488
rect 1211 -1495 1215 -1485
rect 1314 -1472 1318 -1467
rect 940 -1503 1070 -1499
rect 1162 -1500 1203 -1495
rect 1211 -1500 1293 -1495
rect 1162 -1503 1166 -1500
rect 1211 -1503 1215 -1500
rect 975 -1504 1070 -1503
rect 1147 -1507 1184 -1503
rect 1147 -1513 1151 -1507
rect 1180 -1513 1184 -1507
rect 865 -1520 892 -1517
rect 819 -1525 860 -1521
rect 804 -1527 811 -1526
rect 312 -1556 468 -1554
rect 312 -1558 508 -1556
rect 387 -1561 508 -1558
rect 103 -1569 182 -1566
rect 460 -1579 508 -1561
rect 583 -1574 587 -1554
rect 610 -1574 614 -1554
rect 743 -1531 811 -1527
rect 743 -1532 809 -1531
rect 629 -1573 656 -1570
rect 583 -1578 624 -1574
rect 460 -1584 575 -1579
rect 602 -1588 606 -1578
rect 123 -1592 177 -1589
rect 123 -1596 126 -1592
rect 130 -1596 143 -1592
rect 147 -1596 153 -1592
rect 157 -1596 170 -1592
rect 174 -1596 177 -1592
rect 123 -1598 177 -1596
rect 131 -1603 135 -1598
rect 158 -1603 162 -1598
rect 294 -1620 390 -1619
rect 294 -1623 480 -1620
rect 294 -1624 508 -1623
rect 383 -1633 508 -1624
rect 139 -1663 143 -1643
rect 166 -1663 170 -1643
rect 472 -1645 508 -1633
rect 594 -1634 598 -1628
rect 619 -1634 624 -1578
rect 629 -1577 632 -1573
rect 636 -1577 649 -1573
rect 653 -1577 656 -1573
rect 629 -1579 656 -1577
rect 637 -1584 641 -1579
rect 645 -1634 649 -1624
rect 743 -1634 748 -1532
rect 838 -1535 842 -1525
rect 830 -1581 834 -1575
rect 855 -1581 860 -1525
rect 865 -1524 868 -1520
rect 872 -1524 885 -1520
rect 889 -1524 892 -1520
rect 865 -1526 892 -1524
rect 873 -1531 877 -1526
rect 1268 -1506 1293 -1500
rect 1268 -1511 1302 -1506
rect 1203 -1529 1207 -1523
rect 1195 -1530 1222 -1529
rect 1139 -1539 1143 -1533
rect 1172 -1539 1176 -1533
rect 1195 -1534 1196 -1530
rect 1200 -1534 1217 -1530
rect 1221 -1534 1222 -1530
rect 1195 -1535 1222 -1534
rect 1131 -1540 1158 -1539
rect 1131 -1544 1132 -1540
rect 1136 -1544 1153 -1540
rect 1157 -1544 1158 -1540
rect 1131 -1545 1158 -1544
rect 1164 -1540 1191 -1539
rect 1164 -1544 1165 -1540
rect 1169 -1544 1186 -1540
rect 1190 -1544 1191 -1540
rect 1164 -1545 1191 -1544
rect 1297 -1555 1302 -1511
rect 1297 -1560 1314 -1555
rect 1322 -1564 1326 -1552
rect 881 -1581 885 -1571
rect 1314 -1568 1326 -1564
rect 1314 -1572 1318 -1568
rect 830 -1585 844 -1581
rect 838 -1586 844 -1585
rect 855 -1586 873 -1581
rect 881 -1582 894 -1581
rect 881 -1586 1080 -1582
rect 594 -1638 608 -1634
rect 602 -1639 608 -1638
rect 619 -1639 637 -1634
rect 645 -1639 748 -1634
rect 764 -1597 830 -1592
rect 472 -1650 594 -1645
rect 602 -1653 606 -1639
rect 645 -1642 649 -1639
rect 185 -1662 212 -1659
rect 139 -1667 180 -1663
rect 67 -1673 131 -1668
rect 158 -1677 162 -1667
rect 150 -1723 154 -1717
rect 175 -1723 180 -1667
rect 185 -1666 188 -1662
rect 192 -1666 205 -1662
rect 209 -1666 212 -1662
rect 185 -1668 212 -1666
rect 193 -1673 197 -1668
rect 285 -1692 475 -1690
rect 285 -1695 510 -1692
rect 386 -1697 510 -1695
rect 201 -1723 205 -1713
rect 468 -1716 510 -1697
rect 637 -1668 641 -1662
rect 629 -1669 656 -1668
rect 629 -1673 630 -1669
rect 634 -1673 651 -1669
rect 655 -1673 656 -1669
rect 629 -1674 656 -1673
rect 594 -1699 598 -1693
rect 586 -1700 613 -1699
rect 586 -1704 587 -1700
rect 591 -1704 608 -1700
rect 612 -1704 613 -1700
rect 586 -1705 613 -1704
rect 764 -1716 769 -1597
rect 838 -1600 842 -1586
rect 881 -1589 885 -1586
rect 888 -1587 1080 -1586
rect 943 -1596 1088 -1587
rect 873 -1615 877 -1609
rect 865 -1616 892 -1615
rect 865 -1620 866 -1616
rect 870 -1620 887 -1616
rect 891 -1620 892 -1616
rect 865 -1621 892 -1620
rect 830 -1646 834 -1640
rect 822 -1647 849 -1646
rect 822 -1651 823 -1647
rect 827 -1651 844 -1647
rect 848 -1651 849 -1647
rect 822 -1652 849 -1651
rect 812 -1661 866 -1658
rect 812 -1665 815 -1661
rect 819 -1665 832 -1661
rect 836 -1665 842 -1661
rect 846 -1665 859 -1661
rect 863 -1665 866 -1661
rect 812 -1667 866 -1665
rect 820 -1672 824 -1667
rect 847 -1672 851 -1667
rect 1059 -1691 1088 -1596
rect 1157 -1597 1184 -1594
rect 1157 -1601 1160 -1597
rect 1164 -1601 1177 -1597
rect 1181 -1601 1184 -1597
rect 1157 -1603 1184 -1601
rect 1165 -1608 1169 -1603
rect 1355 -1598 1382 -1595
rect 1355 -1602 1358 -1598
rect 1362 -1602 1375 -1598
rect 1379 -1602 1382 -1598
rect 1355 -1604 1382 -1602
rect 1363 -1609 1367 -1604
rect 1059 -1696 1165 -1691
rect 1173 -1700 1177 -1688
rect 468 -1721 769 -1716
rect 150 -1727 164 -1723
rect 158 -1728 164 -1727
rect 175 -1728 193 -1723
rect 201 -1728 316 -1723
rect 321 -1728 354 -1723
rect 29 -1739 150 -1734
rect -495 -1746 -492 -1742
rect -488 -1746 -470 -1742
rect -466 -1746 -440 -1742
rect -436 -1746 -418 -1742
rect -414 -1746 -388 -1742
rect -384 -1746 -366 -1742
rect -362 -1746 -336 -1742
rect -332 -1746 -314 -1742
rect -310 -1746 -307 -1742
rect -495 -1748 -307 -1746
rect -284 -1746 -280 -1740
rect -252 -1746 -248 -1740
rect 158 -1742 162 -1728
rect 201 -1731 205 -1728
rect -485 -1754 -481 -1748
rect -433 -1754 -429 -1748
rect -381 -1754 -377 -1748
rect -329 -1754 -325 -1748
rect -508 -1803 -485 -1798
rect -508 -1869 -503 -1803
rect -477 -1807 -473 -1794
rect -485 -1811 -473 -1807
rect -455 -1803 -433 -1798
rect -485 -1816 -481 -1811
rect -490 -1865 -485 -1860
rect -477 -1869 -473 -1856
rect -455 -1869 -450 -1803
rect -425 -1807 -421 -1794
rect -373 -1798 -369 -1794
rect -321 -1798 -317 -1794
rect -276 -1798 -272 -1786
rect -244 -1798 -240 -1786
rect 828 -1732 832 -1712
rect 855 -1732 859 -1712
rect 1165 -1704 1177 -1700
rect 1260 -1663 1299 -1658
rect 1322 -1659 1326 -1652
rect 1371 -1659 1375 -1649
rect 1260 -1664 1291 -1663
rect 1322 -1664 1363 -1659
rect 1371 -1664 1443 -1659
rect 1165 -1708 1169 -1704
rect 874 -1731 901 -1728
rect 828 -1736 869 -1732
rect 813 -1738 820 -1737
rect 749 -1742 820 -1738
rect 749 -1743 816 -1742
rect 193 -1757 197 -1751
rect 185 -1758 212 -1757
rect 185 -1762 186 -1758
rect 190 -1762 207 -1758
rect 211 -1762 212 -1758
rect 185 -1763 212 -1762
rect 563 -1774 617 -1771
rect 563 -1778 566 -1774
rect 570 -1778 583 -1774
rect 587 -1778 593 -1774
rect 597 -1778 610 -1774
rect 614 -1778 617 -1774
rect 563 -1780 617 -1778
rect 150 -1788 154 -1782
rect 571 -1785 575 -1780
rect 598 -1785 602 -1780
rect 142 -1789 169 -1788
rect 142 -1793 143 -1789
rect 147 -1793 164 -1789
rect 168 -1793 169 -1789
rect 142 -1794 169 -1793
rect -433 -1811 -421 -1807
rect -403 -1803 -381 -1798
rect -373 -1803 -329 -1798
rect -321 -1803 -284 -1798
rect -276 -1803 -252 -1798
rect -244 -1803 -230 -1798
rect -433 -1816 -429 -1811
rect -438 -1865 -433 -1860
rect -425 -1869 -421 -1856
rect -403 -1869 -398 -1803
rect -384 -1826 -381 -1821
rect -373 -1830 -369 -1803
rect -381 -1861 -377 -1850
rect -381 -1865 -369 -1861
rect -508 -1874 -485 -1869
rect -477 -1874 -433 -1869
rect -425 -1874 -381 -1869
rect -477 -1877 -473 -1874
rect -425 -1877 -421 -1874
rect -373 -1877 -369 -1865
rect -351 -1869 -346 -1803
rect -332 -1826 -329 -1821
rect -321 -1830 -317 -1803
rect -276 -1806 -272 -1803
rect -244 -1806 -240 -1803
rect -284 -1833 -280 -1826
rect -252 -1833 -248 -1826
rect 267 -1825 466 -1824
rect 267 -1829 506 -1825
rect -294 -1835 -230 -1833
rect 385 -1834 506 -1829
rect -294 -1839 -292 -1835
rect -288 -1839 -268 -1835
rect -264 -1839 -260 -1835
rect -256 -1839 -236 -1835
rect -232 -1839 -230 -1835
rect -294 -1841 -230 -1839
rect 459 -1850 506 -1834
rect 579 -1845 583 -1825
rect 606 -1845 610 -1825
rect 625 -1844 652 -1841
rect 579 -1849 620 -1845
rect -329 -1861 -325 -1850
rect 459 -1855 571 -1850
rect 598 -1859 602 -1849
rect -329 -1865 -317 -1861
rect -351 -1874 -329 -1869
rect -321 -1877 -317 -1865
rect 270 -1895 271 -1890
rect 276 -1891 478 -1890
rect 276 -1895 504 -1891
rect -485 -1905 -481 -1897
rect -433 -1905 -429 -1897
rect -381 -1905 -377 -1897
rect -329 -1905 -325 -1897
rect 386 -1905 504 -1895
rect -495 -1906 -307 -1905
rect -495 -1910 -468 -1906
rect -464 -1910 -416 -1906
rect -412 -1910 -364 -1906
rect -360 -1910 -312 -1906
rect -308 -1910 -307 -1906
rect -495 -1911 -307 -1910
rect 470 -1916 504 -1905
rect 590 -1905 594 -1899
rect 615 -1905 620 -1849
rect 625 -1848 628 -1844
rect 632 -1848 645 -1844
rect 649 -1848 652 -1844
rect 625 -1850 652 -1848
rect 633 -1855 637 -1850
rect 641 -1905 645 -1895
rect 749 -1905 754 -1743
rect 847 -1746 851 -1736
rect 839 -1792 843 -1786
rect 864 -1792 869 -1736
rect 874 -1735 877 -1731
rect 881 -1735 894 -1731
rect 898 -1735 901 -1731
rect 874 -1737 901 -1735
rect 882 -1742 886 -1737
rect 890 -1792 894 -1782
rect 1206 -1734 1233 -1731
rect 1206 -1738 1209 -1734
rect 1213 -1738 1226 -1734
rect 1230 -1738 1233 -1734
rect 1206 -1740 1233 -1738
rect 1214 -1745 1218 -1740
rect 839 -1796 853 -1792
rect 847 -1797 853 -1796
rect 864 -1797 882 -1792
rect 890 -1797 928 -1792
rect 1063 -1795 1150 -1794
rect 813 -1804 839 -1803
rect 590 -1909 604 -1905
rect 598 -1910 604 -1909
rect 615 -1910 633 -1905
rect 641 -1910 754 -1905
rect 788 -1808 839 -1804
rect 788 -1809 829 -1808
rect -502 -1924 -495 -1919
rect -490 -1924 -443 -1919
rect -438 -1924 -389 -1919
rect -384 -1924 -337 -1919
rect 470 -1921 590 -1916
rect 470 -1922 504 -1921
rect 598 -1924 602 -1910
rect 641 -1913 645 -1910
rect 633 -1939 637 -1933
rect 625 -1940 652 -1939
rect 625 -1944 626 -1940
rect 630 -1944 647 -1940
rect 651 -1944 652 -1940
rect 625 -1945 652 -1944
rect 590 -1970 594 -1964
rect 582 -1971 609 -1970
rect 582 -1975 583 -1971
rect 587 -1975 604 -1971
rect 608 -1975 609 -1971
rect 582 -1976 609 -1975
rect 551 -2023 605 -2020
rect 551 -2027 554 -2023
rect 558 -2027 571 -2023
rect 575 -2027 581 -2023
rect 585 -2027 598 -2023
rect 602 -2027 605 -2023
rect 551 -2029 605 -2027
rect 559 -2034 563 -2029
rect 586 -2034 590 -2029
rect 306 -2078 307 -2073
rect 312 -2076 471 -2073
rect 312 -2078 507 -2076
rect 384 -2085 507 -2078
rect 462 -2099 507 -2085
rect 567 -2094 571 -2074
rect 594 -2094 598 -2074
rect 613 -2093 640 -2090
rect 567 -2098 608 -2094
rect -278 -2104 -214 -2101
rect 462 -2104 559 -2099
rect -278 -2108 -275 -2104
rect -271 -2108 -253 -2104
rect -249 -2108 -243 -2104
rect -239 -2108 -221 -2104
rect -217 -2108 -214 -2104
rect 586 -2108 590 -2098
rect -479 -2112 -291 -2109
rect -278 -2110 -214 -2108
rect -479 -2116 -476 -2112
rect -472 -2116 -454 -2112
rect -450 -2116 -424 -2112
rect -420 -2116 -402 -2112
rect -398 -2116 -372 -2112
rect -368 -2116 -350 -2112
rect -346 -2116 -320 -2112
rect -316 -2116 -298 -2112
rect -294 -2116 -291 -2112
rect -479 -2118 -291 -2116
rect -268 -2116 -264 -2110
rect -236 -2116 -232 -2110
rect -469 -2124 -465 -2118
rect -417 -2124 -413 -2118
rect -365 -2124 -361 -2118
rect -313 -2124 -309 -2118
rect 294 -2144 511 -2139
rect 384 -2152 511 -2144
rect -492 -2173 -469 -2168
rect -492 -2239 -487 -2173
rect -461 -2177 -457 -2164
rect -469 -2181 -457 -2177
rect -439 -2173 -417 -2168
rect -469 -2186 -465 -2181
rect -474 -2235 -469 -2230
rect -461 -2239 -457 -2226
rect -439 -2239 -434 -2173
rect -409 -2177 -405 -2164
rect -357 -2168 -353 -2164
rect -305 -2168 -301 -2164
rect -260 -2168 -256 -2156
rect -228 -2168 -224 -2156
rect 475 -2165 511 -2152
rect 578 -2154 582 -2148
rect 603 -2154 608 -2098
rect 613 -2097 616 -2093
rect 620 -2097 633 -2093
rect 637 -2097 640 -2093
rect 613 -2099 640 -2097
rect 621 -2104 625 -2099
rect 629 -2154 633 -2144
rect 788 -2154 793 -1809
rect 847 -1811 851 -1797
rect 890 -1800 894 -1797
rect 882 -1826 886 -1820
rect 874 -1827 901 -1826
rect 874 -1831 875 -1827
rect 879 -1831 896 -1827
rect 900 -1831 901 -1827
rect 874 -1832 901 -1831
rect 923 -1844 928 -1797
rect 1060 -1799 1150 -1795
rect 1173 -1795 1177 -1788
rect 1222 -1795 1226 -1785
rect 1260 -1795 1288 -1664
rect 1322 -1667 1326 -1664
rect 1371 -1667 1375 -1664
rect 1307 -1671 1344 -1667
rect 1307 -1677 1311 -1671
rect 1340 -1677 1344 -1671
rect 1363 -1693 1367 -1687
rect 1355 -1694 1382 -1693
rect 1299 -1703 1303 -1697
rect 1332 -1703 1336 -1697
rect 1355 -1698 1356 -1694
rect 1360 -1698 1377 -1694
rect 1381 -1698 1382 -1694
rect 1355 -1699 1382 -1698
rect 1291 -1704 1318 -1703
rect 1291 -1708 1292 -1704
rect 1296 -1708 1313 -1704
rect 1317 -1708 1318 -1704
rect 1291 -1709 1318 -1708
rect 1324 -1704 1351 -1703
rect 1324 -1708 1325 -1704
rect 1329 -1708 1346 -1704
rect 1350 -1708 1351 -1704
rect 1324 -1709 1351 -1708
rect 1421 -1773 1443 -1664
rect 2102 -1743 2166 -1740
rect 2102 -1747 2105 -1743
rect 2109 -1747 2127 -1743
rect 2131 -1747 2137 -1743
rect 2141 -1747 2159 -1743
rect 2163 -1747 2166 -1743
rect 1901 -1751 2089 -1748
rect 2102 -1749 2166 -1747
rect 1584 -1757 1611 -1754
rect 1901 -1755 1904 -1751
rect 1908 -1755 1926 -1751
rect 1930 -1755 1956 -1751
rect 1960 -1755 1978 -1751
rect 1982 -1755 2008 -1751
rect 2012 -1755 2030 -1751
rect 2034 -1755 2060 -1751
rect 2064 -1755 2082 -1751
rect 2086 -1755 2089 -1751
rect 1901 -1757 2089 -1755
rect 2112 -1755 2116 -1749
rect 2144 -1755 2148 -1749
rect 1584 -1761 1587 -1757
rect 1591 -1761 1604 -1757
rect 1608 -1761 1611 -1757
rect 1584 -1763 1611 -1761
rect 1911 -1763 1915 -1757
rect 1963 -1763 1967 -1757
rect 2015 -1763 2019 -1757
rect 2067 -1763 2071 -1757
rect 1592 -1768 1596 -1763
rect 1421 -1776 1451 -1773
rect 1481 -1776 1486 -1774
rect 1421 -1778 1486 -1776
rect 1446 -1781 1486 -1778
rect 1060 -1835 1076 -1799
rect 1173 -1800 1214 -1795
rect 1222 -1800 1288 -1795
rect 1446 -1785 1452 -1784
rect 1446 -1789 1447 -1785
rect 1451 -1789 1452 -1785
rect 1446 -1792 1452 -1789
rect 1481 -1792 1486 -1781
rect 1541 -1787 1550 -1784
rect 1541 -1791 1543 -1787
rect 1547 -1791 1550 -1787
rect 1564 -1791 1577 -1788
rect 1541 -1792 1550 -1791
rect 1446 -1796 1458 -1792
rect 1173 -1803 1177 -1800
rect 1222 -1803 1226 -1800
rect 1158 -1807 1195 -1803
rect 1158 -1813 1162 -1807
rect 1191 -1813 1195 -1807
rect 1446 -1806 1452 -1796
rect 1536 -1796 1550 -1792
rect 1478 -1804 1496 -1800
rect 1541 -1804 1550 -1796
rect 1446 -1810 1447 -1806
rect 1451 -1810 1452 -1806
rect 1446 -1811 1452 -1810
rect 1481 -1814 1486 -1804
rect 1541 -1808 1543 -1804
rect 1547 -1808 1550 -1804
rect 1541 -1811 1550 -1808
rect 1556 -1814 1560 -1811
rect 1510 -1818 1560 -1814
rect 1510 -1823 1514 -1818
rect 1214 -1829 1218 -1823
rect 1433 -1824 1514 -1823
rect 1564 -1824 1568 -1811
rect 1571 -1818 1577 -1791
rect 1600 -1818 1604 -1808
rect 1888 -1812 1911 -1807
rect 1571 -1823 1592 -1818
rect 1600 -1823 1611 -1818
rect 1424 -1828 1514 -1824
rect 1206 -1830 1233 -1829
rect 946 -1844 1078 -1835
rect 1150 -1839 1154 -1833
rect 1183 -1839 1187 -1833
rect 1206 -1834 1207 -1830
rect 1211 -1834 1228 -1830
rect 1232 -1834 1233 -1830
rect 1206 -1835 1233 -1834
rect 923 -1849 1078 -1844
rect 1142 -1840 1169 -1839
rect 1142 -1844 1143 -1840
rect 1147 -1844 1164 -1840
rect 1168 -1844 1169 -1840
rect 1142 -1845 1169 -1844
rect 1175 -1840 1202 -1839
rect 1175 -1844 1176 -1840
rect 1180 -1844 1197 -1840
rect 1201 -1844 1202 -1840
rect 1175 -1845 1202 -1844
rect 839 -1857 843 -1851
rect 946 -1852 1078 -1849
rect 831 -1858 858 -1857
rect 831 -1862 832 -1858
rect 836 -1862 853 -1858
rect 857 -1862 858 -1858
rect 831 -1863 858 -1862
rect 1050 -1925 1271 -1924
rect 1050 -1929 1293 -1925
rect 1050 -1973 1083 -1929
rect 1264 -1935 1293 -1929
rect 1424 -1935 1441 -1828
rect 1446 -1836 1452 -1835
rect 1446 -1840 1447 -1836
rect 1451 -1840 1452 -1836
rect 1446 -1843 1452 -1840
rect 1481 -1843 1486 -1828
rect 1541 -1838 1550 -1835
rect 1541 -1842 1543 -1838
rect 1547 -1842 1550 -1838
rect 1541 -1843 1550 -1842
rect 1446 -1847 1458 -1843
rect 1446 -1857 1452 -1847
rect 1536 -1847 1550 -1843
rect 1478 -1855 1496 -1851
rect 1541 -1855 1550 -1847
rect 1446 -1861 1447 -1857
rect 1451 -1861 1452 -1857
rect 1446 -1862 1452 -1861
rect 1481 -1875 1486 -1855
rect 1541 -1859 1543 -1855
rect 1547 -1859 1550 -1855
rect 1541 -1862 1550 -1859
rect 1600 -1826 1604 -1823
rect 1556 -1875 1560 -1844
rect 1592 -1852 1596 -1846
rect 1584 -1853 1611 -1852
rect 1584 -1857 1585 -1853
rect 1589 -1857 1606 -1853
rect 1610 -1857 1611 -1853
rect 1584 -1858 1611 -1857
rect 1481 -1878 1560 -1875
rect 1888 -1878 1893 -1812
rect 1919 -1816 1923 -1803
rect 1911 -1820 1923 -1816
rect 1941 -1812 1963 -1807
rect 1911 -1825 1915 -1820
rect 1906 -1874 1911 -1869
rect 1919 -1878 1923 -1865
rect 1941 -1878 1946 -1812
rect 1971 -1816 1975 -1803
rect 2023 -1807 2027 -1803
rect 2075 -1807 2079 -1803
rect 2120 -1807 2124 -1795
rect 2152 -1807 2156 -1795
rect 1963 -1820 1975 -1816
rect 1993 -1812 2015 -1807
rect 2023 -1812 2067 -1807
rect 2075 -1812 2112 -1807
rect 2120 -1812 2144 -1807
rect 2152 -1812 2166 -1807
rect 1963 -1825 1967 -1820
rect 1958 -1874 1963 -1869
rect 1971 -1878 1975 -1865
rect 1993 -1878 1998 -1812
rect 2012 -1835 2015 -1830
rect 2023 -1839 2027 -1812
rect 2015 -1870 2019 -1859
rect 2015 -1874 2027 -1870
rect 1888 -1883 1911 -1878
rect 1919 -1883 1963 -1878
rect 1971 -1883 2015 -1878
rect 1919 -1886 1923 -1883
rect 1971 -1886 1975 -1883
rect 2023 -1886 2027 -1874
rect 2045 -1878 2050 -1812
rect 2064 -1835 2067 -1830
rect 2075 -1839 2079 -1812
rect 2120 -1815 2124 -1812
rect 2152 -1815 2156 -1812
rect 2112 -1842 2116 -1835
rect 2144 -1842 2148 -1835
rect 2102 -1844 2166 -1842
rect 2102 -1848 2104 -1844
rect 2108 -1848 2128 -1844
rect 2132 -1848 2136 -1844
rect 2140 -1848 2160 -1844
rect 2164 -1848 2166 -1844
rect 2102 -1850 2166 -1848
rect 2067 -1870 2071 -1859
rect 2067 -1874 2079 -1870
rect 2045 -1883 2067 -1878
rect 2075 -1886 2079 -1874
rect 1911 -1914 1915 -1906
rect 1963 -1914 1967 -1906
rect 2015 -1914 2019 -1906
rect 2067 -1914 2071 -1906
rect 1901 -1915 2089 -1914
rect 1901 -1919 1928 -1915
rect 1932 -1919 1980 -1915
rect 1984 -1919 2032 -1915
rect 2036 -1919 2084 -1915
rect 2088 -1919 2089 -1915
rect 1901 -1920 2089 -1919
rect 1894 -1933 1901 -1928
rect 1906 -1933 1953 -1928
rect 1958 -1933 2007 -1928
rect 2012 -1933 2059 -1928
rect 1264 -1939 1441 -1935
rect 1264 -1940 1440 -1939
rect 945 -1974 1083 -1973
rect 578 -2158 592 -2154
rect 586 -2159 592 -2158
rect 603 -2159 621 -2154
rect 629 -2159 793 -2154
rect 816 -1979 1083 -1974
rect -417 -2181 -405 -2177
rect -387 -2173 -365 -2168
rect -357 -2173 -313 -2168
rect -305 -2173 -268 -2168
rect -260 -2173 -236 -2168
rect -228 -2173 -214 -2168
rect 475 -2170 578 -2165
rect 475 -2172 511 -2170
rect 586 -2173 590 -2159
rect 629 -2162 633 -2159
rect -417 -2186 -413 -2181
rect -422 -2235 -417 -2230
rect -409 -2239 -405 -2226
rect -387 -2239 -382 -2173
rect -368 -2196 -365 -2191
rect -357 -2200 -353 -2173
rect -365 -2231 -361 -2220
rect -365 -2235 -353 -2231
rect -492 -2244 -469 -2239
rect -461 -2244 -417 -2239
rect -409 -2244 -365 -2239
rect -461 -2247 -457 -2244
rect -409 -2247 -405 -2244
rect -357 -2247 -353 -2235
rect -335 -2239 -330 -2173
rect -316 -2196 -313 -2191
rect -305 -2200 -301 -2173
rect -260 -2176 -256 -2173
rect -228 -2176 -224 -2173
rect -268 -2203 -264 -2196
rect -236 -2203 -232 -2196
rect -278 -2205 -214 -2203
rect -278 -2209 -276 -2205
rect -272 -2209 -252 -2205
rect -248 -2209 -244 -2205
rect -240 -2209 -220 -2205
rect -216 -2209 -214 -2205
rect -278 -2211 -214 -2209
rect 621 -2188 625 -2182
rect 613 -2189 640 -2188
rect 613 -2193 614 -2189
rect 618 -2193 635 -2189
rect 639 -2193 640 -2189
rect 613 -2194 640 -2193
rect 578 -2219 582 -2213
rect 570 -2220 597 -2219
rect -313 -2231 -309 -2220
rect 570 -2224 571 -2220
rect 575 -2224 592 -2220
rect 596 -2224 597 -2220
rect 570 -2225 597 -2224
rect -313 -2235 -301 -2231
rect 323 -2233 325 -2228
rect 330 -2229 475 -2228
rect 330 -2233 508 -2229
rect -335 -2244 -313 -2239
rect -305 -2247 -301 -2235
rect 383 -2244 508 -2233
rect 464 -2254 508 -2244
rect 816 -2254 821 -1979
rect 945 -1982 1083 -1979
rect 1050 -1985 1083 -1982
rect 464 -2259 821 -2254
rect -469 -2275 -465 -2267
rect -417 -2275 -413 -2267
rect -365 -2275 -361 -2267
rect -313 -2275 -309 -2267
rect -479 -2276 -291 -2275
rect -479 -2280 -452 -2276
rect -448 -2280 -400 -2276
rect -396 -2280 -348 -2276
rect -344 -2280 -296 -2276
rect -292 -2280 -291 -2276
rect -479 -2281 -291 -2280
rect -486 -2294 -479 -2289
rect -474 -2294 -427 -2289
rect -422 -2294 -373 -2289
rect -368 -2294 -321 -2289
rect 599 -2297 1307 -2292
rect 599 -2305 616 -2297
rect 486 -2310 619 -2305
rect 203 -2323 230 -2320
rect 203 -2327 206 -2323
rect 210 -2327 223 -2323
rect 227 -2327 230 -2323
rect 203 -2329 230 -2327
rect 211 -2334 215 -2329
rect 100 -2342 105 -2340
rect -62 -2347 -29 -2342
rect -24 -2347 105 -2342
rect 65 -2351 71 -2350
rect 65 -2355 66 -2351
rect 70 -2355 71 -2351
rect 65 -2358 71 -2355
rect 100 -2358 105 -2347
rect 160 -2353 169 -2350
rect 160 -2357 162 -2353
rect 166 -2357 169 -2353
rect 183 -2357 196 -2354
rect 160 -2358 169 -2357
rect 65 -2362 77 -2358
rect 65 -2372 71 -2362
rect 155 -2362 169 -2358
rect 97 -2370 115 -2366
rect 160 -2370 169 -2362
rect 65 -2376 66 -2372
rect 70 -2376 71 -2372
rect 65 -2377 71 -2376
rect 100 -2380 105 -2370
rect 160 -2374 162 -2370
rect 166 -2374 169 -2370
rect 160 -2377 169 -2374
rect 175 -2380 179 -2377
rect 129 -2384 179 -2380
rect 129 -2389 133 -2384
rect -59 -2394 133 -2389
rect 183 -2390 187 -2377
rect 190 -2384 196 -2357
rect 219 -2384 223 -2374
rect 190 -2389 211 -2384
rect 219 -2389 325 -2384
rect 330 -2389 350 -2384
rect -269 -2533 -205 -2530
rect -269 -2537 -266 -2533
rect -262 -2537 -244 -2533
rect -240 -2537 -234 -2533
rect -230 -2537 -212 -2533
rect -208 -2537 -205 -2533
rect -470 -2541 -282 -2538
rect -269 -2539 -205 -2537
rect -470 -2545 -467 -2541
rect -463 -2545 -445 -2541
rect -441 -2545 -415 -2541
rect -411 -2545 -393 -2541
rect -389 -2545 -363 -2541
rect -359 -2545 -341 -2541
rect -337 -2545 -311 -2541
rect -307 -2545 -289 -2541
rect -285 -2545 -282 -2541
rect -470 -2547 -282 -2545
rect -259 -2545 -255 -2539
rect -227 -2545 -223 -2539
rect -460 -2553 -456 -2547
rect -408 -2553 -404 -2547
rect -356 -2553 -352 -2547
rect -304 -2553 -300 -2547
rect -483 -2602 -460 -2597
rect -483 -2668 -478 -2602
rect -452 -2606 -448 -2593
rect -460 -2610 -448 -2606
rect -430 -2602 -408 -2597
rect -460 -2615 -456 -2610
rect -465 -2664 -460 -2659
rect -452 -2668 -448 -2655
rect -430 -2668 -425 -2602
rect -400 -2606 -396 -2593
rect -348 -2597 -344 -2593
rect -296 -2597 -292 -2593
rect -251 -2597 -247 -2585
rect -219 -2597 -215 -2585
rect -408 -2610 -396 -2606
rect -378 -2602 -356 -2597
rect -348 -2602 -304 -2597
rect -296 -2602 -259 -2597
rect -251 -2602 -227 -2597
rect -219 -2602 -205 -2597
rect -408 -2615 -404 -2610
rect -413 -2664 -408 -2659
rect -400 -2668 -396 -2655
rect -378 -2668 -373 -2602
rect -359 -2625 -356 -2620
rect -348 -2629 -344 -2602
rect -356 -2660 -352 -2649
rect -356 -2664 -344 -2660
rect -483 -2673 -460 -2668
rect -452 -2673 -408 -2668
rect -400 -2673 -356 -2668
rect -452 -2676 -448 -2673
rect -400 -2676 -396 -2673
rect -348 -2676 -344 -2664
rect -326 -2668 -321 -2602
rect -307 -2625 -304 -2620
rect -296 -2629 -292 -2602
rect -251 -2605 -247 -2602
rect -219 -2605 -215 -2602
rect 26 -2609 31 -2394
rect 65 -2402 71 -2401
rect 65 -2406 66 -2402
rect 70 -2406 71 -2402
rect 65 -2409 71 -2406
rect 100 -2409 105 -2394
rect 160 -2404 169 -2401
rect 160 -2408 162 -2404
rect 166 -2408 169 -2404
rect 160 -2409 169 -2408
rect 65 -2413 77 -2409
rect 65 -2423 71 -2413
rect 155 -2413 169 -2409
rect 97 -2421 115 -2417
rect 160 -2421 169 -2413
rect 65 -2427 66 -2423
rect 70 -2427 71 -2423
rect 65 -2428 71 -2427
rect 100 -2441 105 -2421
rect 160 -2425 162 -2421
rect 166 -2425 169 -2421
rect 160 -2428 169 -2425
rect 219 -2392 223 -2389
rect 175 -2441 179 -2410
rect 211 -2418 215 -2412
rect 203 -2419 230 -2418
rect 203 -2423 204 -2419
rect 208 -2423 225 -2419
rect 229 -2423 230 -2419
rect 203 -2424 230 -2423
rect 100 -2444 179 -2441
rect 120 -2467 174 -2464
rect 120 -2471 123 -2467
rect 127 -2471 140 -2467
rect 144 -2471 150 -2467
rect 154 -2471 167 -2467
rect 171 -2471 174 -2467
rect 120 -2473 174 -2471
rect 128 -2478 132 -2473
rect 155 -2478 159 -2473
rect 136 -2538 140 -2518
rect 163 -2538 167 -2518
rect 182 -2537 209 -2534
rect 136 -2542 177 -2538
rect 64 -2548 128 -2543
rect 155 -2552 159 -2542
rect 147 -2598 151 -2592
rect 172 -2598 177 -2542
rect 182 -2541 185 -2537
rect 189 -2541 202 -2537
rect 206 -2541 209 -2537
rect 182 -2543 209 -2541
rect 190 -2548 194 -2543
rect 198 -2598 202 -2588
rect 486 -2598 491 -2310
rect 599 -2311 616 -2310
rect 909 -2328 1277 -2323
rect 690 -2333 744 -2330
rect 690 -2337 693 -2333
rect 697 -2337 710 -2333
rect 714 -2337 720 -2333
rect 724 -2337 737 -2333
rect 741 -2337 744 -2333
rect 690 -2339 744 -2337
rect 698 -2344 702 -2339
rect 725 -2344 729 -2339
rect 706 -2404 710 -2384
rect 733 -2404 737 -2384
rect 752 -2403 779 -2400
rect 706 -2408 747 -2404
rect 599 -2414 698 -2409
rect 601 -2422 618 -2414
rect 725 -2418 729 -2408
rect 147 -2602 161 -2598
rect 155 -2603 161 -2602
rect 172 -2603 190 -2598
rect 198 -2603 491 -2598
rect 500 -2427 619 -2422
rect 26 -2614 147 -2609
rect 155 -2617 159 -2603
rect 198 -2606 202 -2603
rect -259 -2632 -255 -2625
rect -227 -2632 -223 -2625
rect -269 -2634 -205 -2632
rect -269 -2638 -267 -2634
rect -263 -2638 -243 -2634
rect -239 -2638 -235 -2634
rect -231 -2638 -211 -2634
rect -207 -2638 -205 -2634
rect -269 -2640 -205 -2638
rect -304 -2660 -300 -2649
rect 500 -2615 505 -2427
rect 601 -2428 618 -2427
rect 717 -2464 721 -2458
rect 742 -2464 747 -2408
rect 752 -2407 755 -2403
rect 759 -2407 772 -2403
rect 776 -2407 779 -2403
rect 752 -2409 779 -2407
rect 760 -2414 764 -2409
rect 768 -2464 772 -2454
rect 909 -2464 914 -2328
rect 1025 -2385 1079 -2382
rect 1025 -2389 1028 -2385
rect 1032 -2389 1045 -2385
rect 1049 -2389 1055 -2385
rect 1059 -2389 1072 -2385
rect 1076 -2389 1079 -2385
rect 1025 -2391 1079 -2389
rect 1033 -2396 1037 -2391
rect 1060 -2396 1064 -2391
rect 1041 -2456 1045 -2436
rect 1068 -2456 1072 -2436
rect 1087 -2455 1114 -2452
rect 1041 -2460 1082 -2456
rect 717 -2468 731 -2464
rect 725 -2469 731 -2468
rect 742 -2469 760 -2464
rect 768 -2469 914 -2464
rect 1022 -2466 1033 -2461
rect 599 -2480 717 -2475
rect 600 -2488 617 -2480
rect 725 -2483 729 -2469
rect 768 -2472 772 -2469
rect 315 -2620 316 -2615
rect 321 -2620 505 -2615
rect 513 -2493 619 -2488
rect 513 -2624 518 -2493
rect 1022 -2479 1030 -2466
rect 1060 -2470 1064 -2460
rect 961 -2481 1030 -2479
rect 914 -2486 1030 -2481
rect 760 -2498 764 -2492
rect 752 -2499 779 -2498
rect 752 -2503 753 -2499
rect 757 -2503 774 -2499
rect 778 -2503 779 -2499
rect 752 -2504 779 -2503
rect 717 -2529 721 -2523
rect 709 -2530 736 -2529
rect 709 -2534 710 -2530
rect 714 -2534 731 -2530
rect 735 -2534 736 -2530
rect 709 -2535 736 -2534
rect 691 -2616 745 -2613
rect 691 -2620 694 -2616
rect 698 -2620 711 -2616
rect 715 -2620 721 -2616
rect 725 -2620 738 -2616
rect 742 -2620 745 -2616
rect 691 -2622 745 -2620
rect 190 -2632 194 -2626
rect 330 -2629 518 -2624
rect 699 -2627 703 -2622
rect 726 -2627 730 -2622
rect 182 -2633 209 -2632
rect 182 -2637 183 -2633
rect 187 -2637 204 -2633
rect 208 -2637 209 -2633
rect 182 -2638 209 -2637
rect -304 -2664 -292 -2660
rect 147 -2663 151 -2657
rect -326 -2673 -304 -2668
rect -296 -2676 -292 -2664
rect 139 -2664 166 -2663
rect 139 -2668 140 -2664
rect 144 -2668 161 -2664
rect 165 -2668 166 -2664
rect 139 -2669 166 -2668
rect 707 -2687 711 -2667
rect 734 -2687 738 -2667
rect 753 -2686 780 -2683
rect 707 -2691 748 -2687
rect -460 -2704 -456 -2696
rect -408 -2704 -404 -2696
rect -356 -2704 -352 -2696
rect -304 -2704 -300 -2696
rect 599 -2697 699 -2692
rect -470 -2705 -282 -2704
rect 601 -2705 617 -2697
rect 726 -2701 730 -2691
rect -470 -2709 -443 -2705
rect -439 -2709 -391 -2705
rect -387 -2709 -339 -2705
rect -335 -2709 -287 -2705
rect -283 -2709 -282 -2705
rect -470 -2710 -282 -2709
rect 324 -2710 325 -2705
rect 330 -2710 619 -2705
rect -477 -2723 -470 -2718
rect -465 -2723 -418 -2718
rect -413 -2723 -364 -2718
rect -359 -2723 -312 -2718
rect 718 -2747 722 -2741
rect 743 -2747 748 -2691
rect 753 -2690 756 -2686
rect 760 -2690 773 -2686
rect 777 -2690 780 -2686
rect 753 -2692 780 -2690
rect 761 -2697 765 -2692
rect 769 -2747 773 -2737
rect 914 -2747 919 -2486
rect 961 -2487 1030 -2486
rect 1052 -2516 1056 -2510
rect 1077 -2516 1082 -2460
rect 1087 -2459 1090 -2455
rect 1094 -2459 1107 -2455
rect 1111 -2459 1114 -2455
rect 1087 -2461 1114 -2459
rect 1095 -2466 1099 -2461
rect 1103 -2516 1107 -2506
rect 1052 -2520 1066 -2516
rect 1060 -2521 1066 -2520
rect 1077 -2521 1095 -2516
rect 1103 -2521 1261 -2516
rect 718 -2751 732 -2747
rect 726 -2752 732 -2751
rect 743 -2752 761 -2747
rect 769 -2752 919 -2747
rect 951 -2532 1052 -2527
rect 599 -2763 718 -2758
rect 600 -2771 618 -2763
rect 726 -2766 730 -2752
rect 769 -2755 773 -2752
rect 306 -2776 307 -2771
rect 312 -2776 619 -2771
rect 600 -2777 618 -2776
rect 761 -2781 765 -2775
rect 753 -2782 780 -2781
rect 753 -2786 754 -2782
rect 758 -2786 775 -2782
rect 779 -2786 780 -2782
rect 753 -2787 780 -2786
rect 718 -2812 722 -2806
rect 710 -2813 737 -2812
rect 710 -2817 711 -2813
rect 715 -2817 732 -2813
rect 736 -2817 737 -2813
rect 710 -2818 737 -2817
rect 951 -2832 956 -2532
rect 1060 -2535 1064 -2521
rect 1103 -2524 1107 -2521
rect 1095 -2550 1099 -2544
rect 1087 -2551 1114 -2550
rect 1087 -2555 1088 -2551
rect 1092 -2555 1109 -2551
rect 1113 -2555 1114 -2551
rect 1087 -2556 1114 -2555
rect 1052 -2581 1056 -2575
rect 1044 -2582 1071 -2581
rect 1044 -2586 1045 -2582
rect 1049 -2586 1066 -2582
rect 1070 -2586 1071 -2582
rect 1044 -2587 1071 -2586
rect 1026 -2668 1080 -2665
rect 1026 -2672 1029 -2668
rect 1033 -2672 1046 -2668
rect 1050 -2672 1056 -2668
rect 1060 -2672 1073 -2668
rect 1077 -2672 1080 -2668
rect 1026 -2674 1080 -2672
rect 1034 -2679 1038 -2674
rect 1061 -2679 1065 -2674
rect 1042 -2739 1046 -2719
rect 1069 -2739 1073 -2719
rect 1088 -2738 1115 -2735
rect 1042 -2743 1083 -2739
rect 599 -2833 956 -2832
rect 597 -2837 956 -2833
rect 962 -2749 1034 -2744
rect 597 -2845 617 -2837
rect 297 -2850 298 -2845
rect 303 -2850 619 -2845
rect 962 -2850 967 -2749
rect 1061 -2753 1065 -2743
rect 1053 -2799 1057 -2793
rect 1078 -2799 1083 -2743
rect 1088 -2742 1091 -2738
rect 1095 -2742 1108 -2738
rect 1112 -2742 1115 -2738
rect 1088 -2744 1115 -2742
rect 1096 -2749 1100 -2744
rect 1104 -2799 1108 -2789
rect 1053 -2803 1067 -2799
rect 1061 -2804 1067 -2803
rect 1078 -2804 1096 -2799
rect 1104 -2804 1244 -2799
rect 795 -2855 967 -2850
rect 979 -2815 1053 -2810
rect 687 -2887 741 -2884
rect 687 -2891 690 -2887
rect 694 -2891 707 -2887
rect 711 -2891 717 -2887
rect 721 -2891 734 -2887
rect 738 -2891 741 -2887
rect 687 -2893 741 -2891
rect 695 -2898 699 -2893
rect 722 -2898 726 -2893
rect 703 -2958 707 -2938
rect 730 -2958 734 -2938
rect 749 -2957 776 -2954
rect 703 -2962 744 -2958
rect 598 -2968 695 -2963
rect 598 -2976 618 -2968
rect 722 -2972 726 -2962
rect 330 -2981 619 -2976
rect 714 -3018 718 -3012
rect 739 -3018 744 -2962
rect 749 -2961 752 -2957
rect 756 -2961 769 -2957
rect 773 -2961 776 -2957
rect 749 -2963 776 -2961
rect 757 -2968 761 -2963
rect 765 -3018 769 -3008
rect 795 -3018 800 -2855
rect 979 -2872 984 -2815
rect 1061 -2818 1065 -2804
rect 1104 -2807 1108 -2804
rect 1096 -2833 1100 -2827
rect 1088 -2834 1115 -2833
rect 1088 -2838 1089 -2834
rect 1093 -2838 1110 -2834
rect 1114 -2838 1115 -2834
rect 1088 -2839 1115 -2838
rect 1053 -2864 1057 -2858
rect 1045 -2865 1072 -2864
rect 1045 -2869 1046 -2865
rect 1050 -2869 1067 -2865
rect 1071 -2869 1072 -2865
rect 1045 -2870 1072 -2869
rect 714 -3022 728 -3018
rect 722 -3023 728 -3022
rect 739 -3023 757 -3018
rect 765 -3023 800 -3018
rect 809 -2877 984 -2872
rect 599 -3034 714 -3029
rect 599 -3042 619 -3034
rect 722 -3037 726 -3023
rect 765 -3026 769 -3023
rect 306 -3047 307 -3042
rect 312 -3047 619 -3042
rect 757 -3052 761 -3046
rect 749 -3053 776 -3052
rect 749 -3057 750 -3053
rect 754 -3057 771 -3053
rect 775 -3057 776 -3053
rect 749 -3058 776 -3057
rect 714 -3083 718 -3077
rect 706 -3084 733 -3083
rect 706 -3088 707 -3084
rect 711 -3088 728 -3084
rect 732 -3088 733 -3084
rect 706 -3089 733 -3088
rect 675 -3136 729 -3133
rect 675 -3140 678 -3136
rect 682 -3140 695 -3136
rect 699 -3140 705 -3136
rect 709 -3140 722 -3136
rect 726 -3140 729 -3136
rect 675 -3142 729 -3140
rect 683 -3147 687 -3142
rect 710 -3147 714 -3142
rect 691 -3207 695 -3187
rect 718 -3207 722 -3187
rect 737 -3206 764 -3203
rect 691 -3211 732 -3207
rect 599 -3217 683 -3212
rect 599 -3225 618 -3217
rect 710 -3221 714 -3211
rect 285 -3230 619 -3225
rect 702 -3267 706 -3261
rect 727 -3267 732 -3211
rect 737 -3210 740 -3206
rect 744 -3210 757 -3206
rect 761 -3210 764 -3206
rect 737 -3212 764 -3210
rect 745 -3217 749 -3212
rect 753 -3267 757 -3257
rect 809 -3267 814 -2877
rect 1239 -2912 1244 -2804
rect 1256 -2809 1261 -2521
rect 1272 -2523 1277 -2328
rect 1302 -2420 1307 -2297
rect 1355 -2326 1382 -2323
rect 1355 -2330 1358 -2326
rect 1362 -2330 1375 -2326
rect 1379 -2330 1382 -2326
rect 1355 -2332 1382 -2330
rect 1363 -2337 1367 -2332
rect 2090 -2350 2117 -2347
rect 2090 -2354 2093 -2350
rect 2097 -2354 2110 -2350
rect 2114 -2354 2117 -2350
rect 2090 -2356 2117 -2354
rect 1302 -2425 1363 -2420
rect 1302 -2426 1307 -2425
rect 1371 -2429 1375 -2417
rect 1363 -2433 1375 -2429
rect 2098 -2361 2102 -2356
rect 1363 -2437 1367 -2433
rect 2632 -2424 2696 -2421
rect 2632 -2428 2635 -2424
rect 2639 -2428 2657 -2424
rect 2661 -2428 2667 -2424
rect 2671 -2428 2689 -2424
rect 2693 -2428 2696 -2424
rect 2431 -2432 2619 -2429
rect 2632 -2430 2696 -2428
rect 2431 -2436 2434 -2432
rect 2438 -2436 2456 -2432
rect 2460 -2436 2486 -2432
rect 2490 -2436 2508 -2432
rect 2512 -2436 2538 -2432
rect 2542 -2436 2560 -2432
rect 2564 -2436 2590 -2432
rect 2594 -2436 2612 -2432
rect 2616 -2436 2619 -2432
rect 2431 -2438 2619 -2436
rect 2642 -2436 2646 -2430
rect 2674 -2436 2678 -2430
rect 2081 -2445 2098 -2444
rect 1919 -2449 2098 -2445
rect 1919 -2450 2083 -2449
rect 1404 -2463 1431 -2460
rect 1404 -2467 1407 -2463
rect 1411 -2467 1424 -2463
rect 1428 -2467 1431 -2463
rect 1404 -2469 1431 -2467
rect 1412 -2474 1416 -2469
rect 1272 -2528 1348 -2523
rect 1371 -2524 1375 -2517
rect 1420 -2524 1424 -2514
rect 1919 -2524 1924 -2450
rect 2106 -2453 2110 -2441
rect 1371 -2529 1412 -2524
rect 1420 -2529 1924 -2524
rect 2098 -2457 2110 -2453
rect 2441 -2444 2445 -2438
rect 2493 -2444 2497 -2438
rect 2545 -2444 2549 -2438
rect 2597 -2444 2601 -2438
rect 2098 -2461 2102 -2457
rect 1371 -2532 1375 -2529
rect 1420 -2532 1424 -2529
rect 1356 -2536 1393 -2532
rect 1356 -2542 1360 -2536
rect 1389 -2542 1393 -2536
rect 2139 -2487 2166 -2484
rect 2139 -2491 2142 -2487
rect 2146 -2491 2159 -2487
rect 2163 -2491 2166 -2487
rect 2139 -2493 2166 -2491
rect 2418 -2493 2441 -2488
rect 2147 -2498 2151 -2493
rect 2074 -2548 2083 -2547
rect 1967 -2552 2083 -2548
rect 2106 -2548 2110 -2541
rect 2155 -2548 2159 -2538
rect 1412 -2558 1416 -2552
rect 1967 -2553 2076 -2552
rect 2106 -2553 2147 -2548
rect 2155 -2553 2188 -2548
rect 1404 -2559 1431 -2558
rect 1348 -2568 1352 -2562
rect 1381 -2568 1385 -2562
rect 1404 -2563 1405 -2559
rect 1409 -2563 1426 -2559
rect 1430 -2563 1431 -2559
rect 1404 -2564 1431 -2563
rect 1340 -2569 1367 -2568
rect 1340 -2573 1341 -2569
rect 1345 -2573 1362 -2569
rect 1366 -2573 1367 -2569
rect 1340 -2574 1367 -2573
rect 1373 -2569 1400 -2568
rect 1373 -2573 1374 -2569
rect 1378 -2573 1395 -2569
rect 1399 -2573 1400 -2569
rect 1373 -2574 1400 -2573
rect 1362 -2715 1389 -2712
rect 1362 -2719 1365 -2715
rect 1369 -2719 1382 -2715
rect 1386 -2719 1389 -2715
rect 1362 -2721 1389 -2719
rect 1370 -2726 1374 -2721
rect 1256 -2814 1370 -2809
rect 1378 -2818 1382 -2806
rect 1370 -2822 1382 -2818
rect 1370 -2826 1374 -2822
rect 1411 -2852 1438 -2849
rect 1411 -2856 1414 -2852
rect 1418 -2856 1431 -2852
rect 1435 -2856 1438 -2852
rect 1411 -2858 1438 -2856
rect 1419 -2863 1423 -2858
rect 1654 -2871 1681 -2868
rect 1654 -2875 1657 -2871
rect 1661 -2875 1674 -2871
rect 1678 -2875 1681 -2871
rect 1654 -2877 1681 -2875
rect 1239 -2917 1355 -2912
rect 1378 -2913 1382 -2906
rect 1427 -2913 1431 -2903
rect 1662 -2882 1666 -2877
rect 1378 -2918 1419 -2913
rect 1427 -2918 1632 -2913
rect 1378 -2921 1382 -2918
rect 1427 -2921 1431 -2918
rect 1363 -2925 1400 -2921
rect 1363 -2931 1367 -2925
rect 1396 -2931 1400 -2925
rect 1419 -2947 1423 -2941
rect 1411 -2948 1438 -2947
rect 1355 -2957 1359 -2951
rect 1388 -2957 1392 -2951
rect 1411 -2952 1412 -2948
rect 1416 -2952 1433 -2948
rect 1437 -2952 1438 -2948
rect 1411 -2953 1438 -2952
rect 1347 -2958 1374 -2957
rect 1347 -2962 1348 -2958
rect 1352 -2962 1369 -2958
rect 1373 -2962 1374 -2958
rect 1347 -2963 1374 -2962
rect 1380 -2958 1407 -2957
rect 1380 -2962 1381 -2958
rect 1385 -2962 1402 -2958
rect 1406 -2962 1407 -2958
rect 1380 -2963 1407 -2962
rect 1627 -2966 1632 -2918
rect 1645 -2966 1662 -2965
rect 1627 -2970 1662 -2966
rect 1627 -2971 1651 -2970
rect 1670 -2974 1674 -2962
rect 1662 -2978 1674 -2974
rect 1662 -2982 1666 -2978
rect 1703 -3008 1730 -3005
rect 1703 -3012 1706 -3008
rect 1710 -3012 1723 -3008
rect 1727 -3012 1730 -3008
rect 1703 -3014 1730 -3012
rect 1711 -3019 1715 -3014
rect 1356 -3070 1410 -3067
rect 1356 -3074 1359 -3070
rect 1363 -3074 1376 -3070
rect 1380 -3074 1386 -3070
rect 1390 -3074 1403 -3070
rect 1407 -3074 1410 -3070
rect 1356 -3076 1410 -3074
rect 1613 -3073 1647 -3068
rect 1670 -3069 1674 -3062
rect 1719 -3069 1723 -3059
rect 1967 -3069 1972 -2553
rect 2106 -2556 2110 -2553
rect 2155 -2556 2159 -2553
rect 2091 -2560 2128 -2556
rect 2091 -2566 2095 -2560
rect 2124 -2566 2128 -2560
rect 2418 -2559 2423 -2493
rect 2449 -2497 2453 -2484
rect 2441 -2501 2453 -2497
rect 2471 -2493 2493 -2488
rect 2441 -2506 2445 -2501
rect 2436 -2555 2441 -2550
rect 2449 -2559 2453 -2546
rect 2471 -2559 2476 -2493
rect 2501 -2497 2505 -2484
rect 2553 -2488 2557 -2484
rect 2605 -2488 2609 -2484
rect 2650 -2488 2654 -2476
rect 2682 -2488 2686 -2476
rect 2493 -2501 2505 -2497
rect 2523 -2493 2545 -2488
rect 2553 -2493 2597 -2488
rect 2605 -2493 2642 -2488
rect 2650 -2493 2674 -2488
rect 2682 -2493 2696 -2488
rect 2493 -2506 2497 -2501
rect 2488 -2555 2493 -2550
rect 2501 -2559 2505 -2546
rect 2523 -2559 2528 -2493
rect 2542 -2516 2545 -2511
rect 2553 -2520 2557 -2493
rect 2545 -2551 2549 -2540
rect 2545 -2555 2557 -2551
rect 2418 -2564 2441 -2559
rect 2449 -2564 2493 -2559
rect 2501 -2564 2545 -2559
rect 2449 -2567 2453 -2564
rect 2501 -2567 2505 -2564
rect 2553 -2567 2557 -2555
rect 2575 -2559 2580 -2493
rect 2594 -2516 2597 -2511
rect 2605 -2520 2609 -2493
rect 2650 -2496 2654 -2493
rect 2682 -2496 2686 -2493
rect 2642 -2523 2646 -2516
rect 2674 -2523 2678 -2516
rect 2632 -2525 2696 -2523
rect 2632 -2529 2634 -2525
rect 2638 -2529 2658 -2525
rect 2662 -2529 2666 -2525
rect 2670 -2529 2690 -2525
rect 2694 -2529 2696 -2525
rect 2632 -2531 2696 -2529
rect 2597 -2551 2601 -2540
rect 2597 -2555 2609 -2551
rect 2575 -2564 2597 -2559
rect 2605 -2567 2609 -2555
rect 2147 -2582 2151 -2576
rect 2139 -2583 2166 -2582
rect 2083 -2592 2087 -2586
rect 2116 -2592 2120 -2586
rect 2139 -2587 2140 -2583
rect 2144 -2587 2161 -2583
rect 2165 -2587 2166 -2583
rect 2139 -2588 2166 -2587
rect 2075 -2593 2102 -2592
rect 2075 -2597 2076 -2593
rect 2080 -2597 2097 -2593
rect 2101 -2597 2102 -2593
rect 2075 -2598 2102 -2597
rect 2108 -2593 2135 -2592
rect 2108 -2597 2109 -2593
rect 2113 -2597 2130 -2593
rect 2134 -2597 2135 -2593
rect 2441 -2595 2445 -2587
rect 2493 -2595 2497 -2587
rect 2545 -2595 2549 -2587
rect 2597 -2595 2601 -2587
rect 2108 -2598 2135 -2597
rect 2431 -2596 2619 -2595
rect 2431 -2600 2458 -2596
rect 2462 -2600 2510 -2596
rect 2514 -2600 2562 -2596
rect 2566 -2600 2614 -2596
rect 2618 -2600 2619 -2596
rect 2431 -2601 2619 -2600
rect 2424 -2614 2431 -2609
rect 2436 -2614 2483 -2609
rect 2488 -2614 2537 -2609
rect 2542 -2614 2589 -2609
rect 1364 -3081 1368 -3076
rect 1391 -3081 1395 -3076
rect 1372 -3141 1376 -3121
rect 1399 -3141 1403 -3121
rect 1418 -3140 1445 -3137
rect 702 -3271 716 -3267
rect 710 -3272 716 -3271
rect 727 -3272 745 -3267
rect 753 -3272 814 -3267
rect 819 -3146 1361 -3142
rect 1372 -3145 1413 -3141
rect 819 -3147 1364 -3146
rect 599 -3283 702 -3278
rect 600 -3291 618 -3283
rect 710 -3286 714 -3272
rect 753 -3275 757 -3272
rect 288 -3296 289 -3291
rect 294 -3296 619 -3291
rect 745 -3301 749 -3295
rect 737 -3302 764 -3301
rect 737 -3306 738 -3302
rect 742 -3306 759 -3302
rect 763 -3306 764 -3302
rect 737 -3307 764 -3306
rect 702 -3332 706 -3326
rect 694 -3333 721 -3332
rect 694 -3337 695 -3333
rect 699 -3337 716 -3333
rect 720 -3337 721 -3333
rect 694 -3338 721 -3337
rect 692 -3403 746 -3400
rect 692 -3407 695 -3403
rect 699 -3407 712 -3403
rect 716 -3407 722 -3403
rect 726 -3407 739 -3403
rect 743 -3407 746 -3403
rect 692 -3409 746 -3407
rect 700 -3414 704 -3409
rect 727 -3414 731 -3409
rect 708 -3474 712 -3454
rect 735 -3474 739 -3454
rect 754 -3473 781 -3470
rect 708 -3478 749 -3474
rect 599 -3480 700 -3479
rect 598 -3484 700 -3480
rect 598 -3492 618 -3484
rect 727 -3488 731 -3478
rect 261 -3497 262 -3492
rect 267 -3497 619 -3492
rect 719 -3534 723 -3528
rect 744 -3534 749 -3478
rect 754 -3477 757 -3473
rect 761 -3477 774 -3473
rect 778 -3477 781 -3473
rect 754 -3479 781 -3477
rect 762 -3484 766 -3479
rect 770 -3534 774 -3524
rect 819 -3534 824 -3147
rect 1356 -3151 1364 -3147
rect 1356 -3152 1361 -3151
rect 1391 -3155 1395 -3145
rect 1016 -3202 1070 -3199
rect 1016 -3206 1019 -3202
rect 1023 -3206 1036 -3202
rect 1040 -3206 1046 -3202
rect 1050 -3206 1063 -3202
rect 1067 -3206 1070 -3202
rect 1383 -3201 1387 -3195
rect 1408 -3201 1413 -3145
rect 1418 -3144 1421 -3140
rect 1425 -3144 1438 -3140
rect 1442 -3144 1445 -3140
rect 1418 -3146 1445 -3144
rect 1426 -3151 1430 -3146
rect 1434 -3201 1438 -3191
rect 1613 -3201 1618 -3073
rect 1670 -3074 1711 -3069
rect 1719 -3074 1972 -3069
rect 1670 -3077 1674 -3074
rect 1719 -3077 1723 -3074
rect 1655 -3081 1692 -3077
rect 1655 -3087 1659 -3081
rect 1688 -3087 1692 -3081
rect 1711 -3103 1715 -3097
rect 1703 -3104 1730 -3103
rect 1647 -3113 1651 -3107
rect 1680 -3113 1684 -3107
rect 1703 -3108 1704 -3104
rect 1708 -3108 1725 -3104
rect 1729 -3108 1730 -3104
rect 1703 -3109 1730 -3108
rect 1639 -3114 1666 -3113
rect 1639 -3118 1640 -3114
rect 1644 -3118 1661 -3114
rect 1665 -3118 1666 -3114
rect 1639 -3119 1666 -3118
rect 1672 -3114 1699 -3113
rect 1672 -3118 1673 -3114
rect 1677 -3118 1694 -3114
rect 1698 -3118 1699 -3114
rect 1672 -3119 1699 -3118
rect 1383 -3205 1397 -3201
rect 1016 -3208 1070 -3206
rect 1391 -3206 1397 -3205
rect 1408 -3206 1426 -3201
rect 1434 -3206 1618 -3201
rect 1024 -3213 1028 -3208
rect 1051 -3213 1055 -3208
rect 1032 -3273 1036 -3253
rect 1059 -3273 1063 -3253
rect 1159 -3217 1383 -3212
rect 1078 -3272 1105 -3269
rect 1017 -3278 1022 -3276
rect 1032 -3277 1073 -3273
rect 1017 -3280 1024 -3278
rect 719 -3538 733 -3534
rect 727 -3539 733 -3538
rect 744 -3539 762 -3534
rect 770 -3539 824 -3534
rect 904 -3283 1024 -3280
rect 904 -3285 1022 -3283
rect 599 -3550 719 -3545
rect 600 -3558 618 -3550
rect 727 -3553 731 -3539
rect 770 -3542 774 -3539
rect 270 -3563 271 -3558
rect 276 -3563 619 -3558
rect 600 -3564 618 -3563
rect 762 -3568 766 -3562
rect 754 -3569 781 -3568
rect 754 -3573 755 -3569
rect 759 -3573 776 -3569
rect 780 -3573 781 -3569
rect 754 -3574 781 -3573
rect 719 -3599 723 -3593
rect 711 -3600 738 -3599
rect 711 -3604 712 -3600
rect 716 -3604 733 -3600
rect 737 -3604 738 -3600
rect 711 -3605 738 -3604
rect 680 -3652 734 -3649
rect 680 -3656 683 -3652
rect 687 -3656 700 -3652
rect 704 -3656 710 -3652
rect 714 -3656 727 -3652
rect 731 -3656 734 -3652
rect 680 -3658 734 -3656
rect 688 -3663 692 -3658
rect 715 -3663 719 -3658
rect 696 -3723 700 -3703
rect 723 -3723 727 -3703
rect 742 -3722 769 -3719
rect 696 -3727 737 -3723
rect 599 -3733 688 -3728
rect 599 -3741 617 -3733
rect 715 -3737 719 -3727
rect 288 -3746 289 -3741
rect 294 -3746 619 -3741
rect 707 -3783 711 -3777
rect 732 -3783 737 -3727
rect 742 -3726 745 -3722
rect 749 -3726 762 -3722
rect 766 -3726 769 -3722
rect 742 -3728 769 -3726
rect 750 -3733 754 -3728
rect 758 -3783 762 -3773
rect 904 -3783 909 -3285
rect 1017 -3287 1022 -3285
rect 1051 -3287 1055 -3277
rect 1043 -3333 1047 -3327
rect 1068 -3333 1073 -3277
rect 1078 -3276 1081 -3272
rect 1085 -3276 1098 -3272
rect 1102 -3276 1105 -3272
rect 1078 -3278 1105 -3276
rect 1086 -3283 1090 -3278
rect 1094 -3333 1098 -3323
rect 1159 -3332 1164 -3217
rect 1391 -3220 1395 -3206
rect 1434 -3209 1438 -3206
rect 1426 -3235 1430 -3229
rect 1418 -3236 1445 -3235
rect 1418 -3240 1419 -3236
rect 1423 -3240 1440 -3236
rect 1444 -3240 1445 -3236
rect 1418 -3241 1445 -3240
rect 1383 -3266 1387 -3260
rect 1375 -3267 1402 -3266
rect 1375 -3271 1376 -3267
rect 1380 -3271 1397 -3267
rect 1401 -3271 1402 -3267
rect 1375 -3272 1402 -3271
rect 1104 -3333 1164 -3332
rect 1043 -3337 1057 -3333
rect 1051 -3338 1057 -3337
rect 1068 -3338 1086 -3333
rect 1094 -3337 1164 -3333
rect 1094 -3338 1107 -3337
rect 707 -3787 721 -3783
rect 715 -3788 721 -3787
rect 732 -3788 750 -3783
rect 758 -3788 909 -3783
rect 950 -3349 1043 -3344
rect 599 -3799 707 -3794
rect 600 -3807 619 -3799
rect 715 -3802 719 -3788
rect 758 -3791 762 -3788
rect 306 -3812 307 -3807
rect 312 -3812 619 -3807
rect 600 -3813 619 -3812
rect 750 -3817 754 -3811
rect 742 -3818 769 -3817
rect 742 -3822 743 -3818
rect 747 -3822 764 -3818
rect 768 -3822 769 -3818
rect 742 -3823 769 -3822
rect 707 -3848 711 -3842
rect 699 -3849 726 -3848
rect 699 -3853 700 -3849
rect 704 -3853 721 -3849
rect 725 -3853 726 -3849
rect 699 -3854 726 -3853
rect 950 -3863 955 -3349
rect 1051 -3352 1055 -3338
rect 1094 -3341 1098 -3338
rect 1086 -3367 1090 -3361
rect 1078 -3368 1105 -3367
rect 1078 -3372 1079 -3368
rect 1083 -3372 1100 -3368
rect 1104 -3372 1105 -3368
rect 1078 -3373 1105 -3372
rect 1043 -3398 1047 -3392
rect 1035 -3399 1062 -3398
rect 1035 -3403 1036 -3399
rect 1040 -3403 1057 -3399
rect 1061 -3403 1062 -3399
rect 1035 -3404 1062 -3403
rect 599 -3868 955 -3863
rect 599 -3876 619 -3868
rect 324 -3881 325 -3876
rect 330 -3881 619 -3876
<< m2contact >>
rect 1161 94 1166 99
rect 1213 94 1218 99
rect 1267 133 1272 138
rect 1319 133 1324 138
rect -470 -32 -465 -27
rect 1161 35 1166 40
rect 1213 35 1218 40
rect 1267 35 1272 40
rect 1319 35 1324 40
rect -418 -32 -413 -27
rect -364 7 -359 12
rect -312 7 -307 12
rect 299 26 304 31
rect 308 -22 313 -17
rect -470 -91 -465 -86
rect -418 -91 -413 -86
rect -364 -91 -359 -86
rect -312 -91 -307 -86
rect 14 -176 19 -171
rect 308 -218 313 -213
rect -437 -427 -432 -422
rect -385 -427 -380 -422
rect -331 -388 -326 -383
rect -279 -388 -274 -383
rect 299 -284 304 -279
rect 101 -377 107 -372
rect 317 -432 322 -427
rect -437 -486 -432 -481
rect -385 -486 -380 -481
rect -331 -486 -326 -481
rect -279 -486 -274 -481
rect 326 -461 331 -456
rect 1439 -369 1444 -364
rect 1491 -369 1496 -364
rect 1545 -330 1550 -325
rect 1597 -330 1602 -325
rect 1439 -428 1444 -423
rect 1491 -428 1496 -423
rect 1545 -428 1550 -423
rect 1597 -428 1602 -423
rect 298 -714 303 -709
rect -546 -806 -541 -801
rect 280 -738 285 -733
rect -494 -806 -489 -801
rect -440 -767 -435 -762
rect -388 -767 -383 -762
rect -35 -812 -30 -807
rect 289 -854 294 -849
rect -546 -865 -541 -860
rect -494 -865 -489 -860
rect -440 -865 -435 -860
rect -388 -865 -383 -860
rect 262 -983 267 -978
rect 271 -995 276 -990
rect 52 -1013 58 -1008
rect 298 -1068 303 -1063
rect -470 -1159 -465 -1154
rect -418 -1159 -413 -1154
rect -364 -1120 -359 -1115
rect -312 -1120 -307 -1115
rect 289 -1121 294 -1116
rect 1750 -924 1755 -919
rect 1802 -924 1807 -919
rect 1856 -885 1861 -880
rect 1908 -885 1913 -880
rect 1750 -983 1755 -978
rect 1802 -983 1807 -978
rect 1856 -983 1861 -978
rect 1908 -983 1913 -978
rect 307 -1155 312 -1149
rect 316 -1169 321 -1164
rect -470 -1218 -465 -1213
rect -418 -1218 -413 -1213
rect -364 -1218 -359 -1213
rect -312 -1218 -307 -1213
rect 307 -1275 312 -1270
rect 298 -1341 303 -1336
rect -479 -1487 -474 -1482
rect -427 -1487 -422 -1482
rect -373 -1448 -368 -1443
rect -321 -1448 -316 -1443
rect -26 -1472 -21 -1467
rect 307 -1514 312 -1509
rect -479 -1546 -474 -1541
rect -427 -1546 -422 -1541
rect -373 -1546 -368 -1541
rect -321 -1546 -316 -1541
rect 307 -1558 312 -1553
rect 289 -1624 294 -1619
rect 61 -1673 67 -1668
rect 280 -1695 285 -1690
rect 316 -1728 321 -1723
rect -495 -1865 -490 -1860
rect -443 -1865 -438 -1860
rect -389 -1826 -384 -1821
rect -337 -1826 -332 -1821
rect 262 -1829 267 -1824
rect 271 -1895 276 -1890
rect -495 -1924 -490 -1919
rect -443 -1924 -438 -1919
rect -389 -1924 -384 -1919
rect -337 -1924 -332 -1919
rect 307 -2078 312 -2073
rect 289 -2144 294 -2139
rect -479 -2235 -474 -2230
rect 1901 -1874 1906 -1869
rect 1953 -1874 1958 -1869
rect 2007 -1835 2012 -1830
rect 2059 -1835 2064 -1830
rect 1901 -1933 1906 -1928
rect 1953 -1933 1958 -1928
rect 2007 -1933 2012 -1928
rect 2059 -1933 2064 -1928
rect -427 -2235 -422 -2230
rect -373 -2196 -368 -2191
rect -321 -2196 -316 -2191
rect 325 -2233 330 -2228
rect -479 -2294 -474 -2289
rect -427 -2294 -422 -2289
rect -373 -2294 -368 -2289
rect -321 -2294 -316 -2289
rect -29 -2347 -24 -2342
rect 325 -2389 330 -2384
rect -470 -2664 -465 -2659
rect -418 -2664 -413 -2659
rect -364 -2625 -359 -2620
rect -312 -2625 -307 -2620
rect 58 -2548 64 -2543
rect 316 -2620 321 -2615
rect 325 -2629 330 -2624
rect 325 -2710 330 -2705
rect -470 -2723 -465 -2718
rect -418 -2723 -413 -2718
rect -364 -2723 -359 -2718
rect -312 -2723 -307 -2718
rect 307 -2776 312 -2771
rect 298 -2850 303 -2845
rect 325 -2981 330 -2976
rect 307 -3047 312 -3042
rect 280 -3230 285 -3225
rect 2431 -2555 2436 -2550
rect 2483 -2555 2488 -2550
rect 2537 -2516 2542 -2511
rect 2589 -2516 2594 -2511
rect 2431 -2614 2436 -2609
rect 2483 -2614 2488 -2609
rect 2537 -2614 2542 -2609
rect 2589 -2614 2594 -2609
rect 289 -3296 294 -3291
rect 262 -3497 267 -3492
rect 271 -3563 276 -3558
rect 289 -3746 294 -3741
rect 307 -3812 312 -3807
rect 325 -3881 330 -3876
<< metal2 >>
rect 1161 40 1166 94
rect 1213 40 1218 94
rect 1267 40 1272 133
rect 1319 40 1324 133
rect -470 -86 -465 -32
rect -418 -86 -413 -32
rect -364 -86 -359 7
rect -312 -86 -307 7
rect 14 -372 19 -176
rect 299 -279 304 26
rect 14 -377 101 -372
rect -437 -481 -432 -427
rect -385 -481 -380 -427
rect -331 -481 -326 -388
rect -279 -481 -274 -388
rect 299 -570 304 -284
rect 262 -574 304 -570
rect 308 -213 313 -22
rect -546 -860 -541 -806
rect -494 -860 -489 -806
rect -440 -860 -435 -767
rect -388 -860 -383 -767
rect -35 -1008 -30 -812
rect 262 -978 267 -574
rect 308 -578 313 -218
rect 1439 -423 1444 -369
rect -35 -1013 52 -1008
rect -470 -1213 -465 -1159
rect -418 -1213 -413 -1159
rect -364 -1213 -359 -1120
rect -312 -1213 -307 -1120
rect -479 -1541 -474 -1487
rect -427 -1541 -422 -1487
rect -373 -1541 -368 -1448
rect -321 -1541 -316 -1448
rect -26 -1668 -21 -1472
rect -26 -1673 61 -1668
rect -495 -1919 -490 -1865
rect -443 -1919 -438 -1865
rect -389 -1919 -384 -1826
rect -337 -1919 -332 -1826
rect 262 -1824 267 -983
rect -479 -2289 -474 -2235
rect -427 -2289 -422 -2235
rect -373 -2289 -368 -2196
rect -321 -2289 -316 -2196
rect -29 -2543 -24 -2347
rect -29 -2548 58 -2543
rect -470 -2718 -465 -2664
rect -418 -2718 -413 -2664
rect -364 -2718 -359 -2625
rect -312 -2718 -307 -2625
rect 262 -3492 267 -1829
rect 262 -3885 267 -3497
rect 271 -581 313 -578
rect 1491 -423 1496 -369
rect 1545 -423 1550 -330
rect 1597 -423 1602 -330
rect 271 -990 276 -581
rect 317 -585 322 -432
rect 271 -1890 276 -995
rect 271 -3558 276 -1895
rect 271 -3886 276 -3563
rect 280 -588 322 -585
rect 280 -733 285 -588
rect 326 -592 331 -461
rect 280 -1690 285 -738
rect 280 -3225 285 -1695
rect 280 -3882 285 -3230
rect 289 -597 331 -592
rect 289 -849 294 -597
rect 289 -1116 294 -854
rect 289 -1619 294 -1121
rect 289 -2139 294 -1624
rect 289 -3291 294 -2144
rect 289 -3741 294 -3296
rect 289 -3884 294 -3746
rect 298 -1063 303 -714
rect 1750 -978 1755 -924
rect 1802 -978 1807 -924
rect 1856 -978 1861 -885
rect 1908 -978 1913 -885
rect 298 -1336 303 -1068
rect 298 -2845 303 -1341
rect 298 -3883 303 -2850
rect 307 -1270 312 -1155
rect 307 -1509 312 -1275
rect 307 -1553 312 -1514
rect 307 -2073 312 -1558
rect 307 -2771 312 -2078
rect 307 -3042 312 -2776
rect 307 -3807 312 -3047
rect 307 -3883 312 -3812
rect 316 -1723 321 -1169
rect 316 -2615 321 -1728
rect 1901 -1928 1906 -1874
rect 1953 -1928 1958 -1874
rect 2007 -1928 2012 -1835
rect 2059 -1928 2064 -1835
rect 316 -3884 321 -2620
rect 325 -2228 330 -2223
rect 325 -2384 330 -2233
rect 325 -2624 330 -2389
rect 2431 -2609 2436 -2555
rect 2483 -2609 2488 -2555
rect 2537 -2609 2542 -2516
rect 2589 -2609 2594 -2516
rect 325 -2705 330 -2629
rect 325 -2976 330 -2710
rect 325 -3876 330 -2981
rect 325 -3884 330 -3881
<< labels >>
rlabel metal1 207 -243 207 -243 7 vdd
rlabel metal1 111 -243 111 -243 3 gnd
rlabel metal1 207 -192 207 -192 7 vdd
rlabel metal1 111 -192 111 -192 3 gnd
rlabel metal1 259 -250 259 -250 1 gnd
rlabel metal1 259 -154 259 -154 5 vdd
rlabel metal1 176 -298 176 -298 5 vdd
rlabel metal1 203 -298 203 -298 5 vdd
rlabel metal1 195 -495 195 -495 1 gnd
rlabel metal1 238 -368 238 -368 5 vdd
rlabel metal1 238 -464 238 -464 1 gnd
rlabel metal1 292 -430 292 -430 1 G0
rlabel metal1 287 -216 287 -216 1 P0
rlabel metal1 -14 28 -14 28 1 c0
rlabel metal1 631 -59 631 -59 1 gnd
rlabel metal1 631 37 631 37 5 vdd
rlabel metal1 483 -1 483 -1 3 gnd
rlabel metal1 579 -1 579 -1 7 vdd
rlabel metal1 483 -52 483 -52 3 gnd
rlabel metal1 579 -52 579 -52 7 vdd
rlabel metal1 1127 -350 1127 -350 5 vdd
rlabel metal1 1127 -446 1127 -446 1 gnd
rlabel metal1 979 -388 979 -388 3 gnd
rlabel metal1 1075 -388 1075 -388 7 vdd
rlabel metal1 979 -439 979 -439 3 gnd
rlabel metal1 1075 -439 1075 -439 7 vdd
rlabel metal1 794 -334 794 -334 1 c1
rlabel metal1 774 -370 774 -370 1 gnd
rlabel metal1 774 -274 774 -274 5 vdd
rlabel metal1 743 -380 743 -380 1 gnd
rlabel metal1 710 -380 710 -380 1 gnd
rlabel metal1 725 -137 725 -137 5 vdd
rlabel metal1 480 -170 480 -170 5 vdd
rlabel metal1 507 -170 507 -170 5 vdd
rlabel metal1 499 -367 499 -367 1 gnd
rlabel metal1 542 -240 542 -240 5 vdd
rlabel metal1 542 -336 542 -336 1 gnd
rlabel metal1 167 -1539 167 -1539 7 vdd
rlabel metal1 71 -1539 71 -1539 3 gnd
rlabel metal1 167 -1488 167 -1488 7 vdd
rlabel metal1 71 -1488 71 -1488 3 gnd
rlabel metal1 219 -1546 219 -1546 1 gnd
rlabel metal1 219 -1450 219 -1450 5 vdd
rlabel metal1 136 -1594 136 -1594 5 vdd
rlabel metal1 163 -1594 163 -1594 5 vdd
rlabel metal1 155 -1791 155 -1791 1 gnd
rlabel metal1 198 -1664 198 -1664 5 vdd
rlabel metal1 198 -1760 198 -1760 1 gnd
rlabel metal1 253 -1512 253 -1512 1 P2
rlabel metal1 250 -1726 250 -1726 1 G2
rlabel metal1 158 -879 158 -879 7 vdd
rlabel metal1 62 -879 62 -879 3 gnd
rlabel metal1 158 -828 158 -828 7 vdd
rlabel metal1 62 -828 62 -828 3 gnd
rlabel metal1 210 -886 210 -886 1 gnd
rlabel metal1 210 -790 210 -790 5 vdd
rlabel metal1 127 -934 127 -934 5 vdd
rlabel metal1 154 -934 154 -934 5 vdd
rlabel metal1 146 -1131 146 -1131 1 gnd
rlabel metal1 189 -1004 189 -1004 5 vdd
rlabel metal1 189 -1100 189 -1100 1 gnd
rlabel metal1 244 -852 244 -852 1 P1
rlabel metal1 244 -1066 244 -1066 1 G1
rlabel metal1 164 -2414 164 -2414 7 vdd
rlabel metal1 68 -2414 68 -2414 3 gnd
rlabel metal1 164 -2363 164 -2363 7 vdd
rlabel metal1 68 -2363 68 -2363 3 gnd
rlabel metal1 216 -2421 216 -2421 1 gnd
rlabel metal1 216 -2325 216 -2325 5 vdd
rlabel metal1 133 -2469 133 -2469 5 vdd
rlabel metal1 160 -2469 160 -2469 5 vdd
rlabel metal1 152 -2666 152 -2666 1 gnd
rlabel metal1 195 -2539 195 -2539 5 vdd
rlabel metal1 195 -2635 195 -2635 1 gnd
rlabel metal1 250 -2387 250 -2387 1 P3
rlabel metal1 247 -2601 247 -2601 1 G3
rlabel metal1 1255 -851 1255 -851 1 gnd
rlabel metal1 1255 -755 1255 -755 5 vdd
rlabel metal1 1224 -861 1224 -861 1 gnd
rlabel metal1 1191 -861 1191 -861 1 gnd
rlabel metal1 1206 -618 1206 -618 5 vdd
rlabel metal1 1481 -795 1481 -795 5 vdd
rlabel metal1 1481 -891 1481 -891 1 gnd
rlabel metal1 1333 -833 1333 -833 3 gnd
rlabel metal1 1429 -833 1429 -833 7 vdd
rlabel metal1 1333 -884 1333 -884 3 gnd
rlabel metal1 1429 -884 1429 -884 7 vdd
rlabel metal1 722 -904 722 -904 5 vdd
rlabel metal1 749 -904 749 -904 5 vdd
rlabel metal1 741 -1101 741 -1101 1 gnd
rlabel metal1 784 -974 784 -974 5 vdd
rlabel metal1 784 -1070 784 -1070 1 gnd
rlabel metal1 504 -904 504 -904 5 vdd
rlabel metal1 531 -904 531 -904 5 vdd
rlabel metal1 523 -1101 523 -1101 1 gnd
rlabel metal1 566 -974 566 -974 5 vdd
rlabel metal1 566 -1070 566 -1070 1 gnd
rlabel metal1 581 -659 581 -659 5 vdd
rlabel metal1 608 -659 608 -659 5 vdd
rlabel metal1 600 -856 600 -856 1 gnd
rlabel metal1 643 -729 643 -729 5 vdd
rlabel metal1 643 -825 643 -825 1 gnd
rlabel metal1 980 -626 980 -626 5 vdd
rlabel metal1 965 -869 965 -869 1 gnd
rlabel metal1 998 -869 998 -869 1 gnd
rlabel metal1 1029 -763 1029 -763 5 vdd
rlabel metal1 1029 -859 1029 -859 1 gnd
rlabel metal1 878 -1522 878 -1522 5 vdd
rlabel metal1 835 -1649 835 -1649 1 gnd
rlabel metal1 843 -1452 843 -1452 5 vdd
rlabel metal1 816 -1452 816 -1452 5 vdd
rlabel metal1 887 -1829 887 -1829 1 gnd
rlabel metal1 887 -1733 887 -1733 5 vdd
rlabel metal1 844 -1860 844 -1860 1 gnd
rlabel metal1 852 -1663 852 -1663 5 vdd
rlabel metal1 825 -1663 825 -1663 5 vdd
rlabel metal1 638 -1942 638 -1942 1 gnd
rlabel metal1 638 -1846 638 -1846 5 vdd
rlabel metal1 595 -1973 595 -1973 1 gnd
rlabel metal1 603 -1776 603 -1776 5 vdd
rlabel metal1 576 -1776 576 -1776 5 vdd
rlabel metal1 642 -1671 642 -1671 1 gnd
rlabel metal1 642 -1575 642 -1575 5 vdd
rlabel metal1 599 -1702 599 -1702 1 gnd
rlabel metal1 607 -1505 607 -1505 5 vdd
rlabel metal1 580 -1505 580 -1505 5 vdd
rlabel metal1 641 -1388 641 -1388 1 gnd
rlabel metal1 641 -1292 641 -1292 5 vdd
rlabel metal1 598 -1419 598 -1419 1 gnd
rlabel metal1 606 -1222 606 -1222 5 vdd
rlabel metal1 579 -1222 579 -1222 5 vdd
rlabel metal1 626 -2191 626 -2191 1 gnd
rlabel metal1 626 -2095 626 -2095 5 vdd
rlabel metal1 591 -2025 591 -2025 5 vdd
rlabel metal1 564 -2025 564 -2025 5 vdd
rlabel metal1 583 -2222 583 -2222 1 gnd
rlabel metal1 878 -1618 878 -1618 1 gnd
rlabel metal1 1597 -1759 1597 -1759 5 vdd
rlabel metal1 1597 -1855 1597 -1855 1 gnd
rlabel metal1 1449 -1797 1449 -1797 3 gnd
rlabel metal1 1545 -1797 1545 -1797 7 vdd
rlabel metal1 1449 -1848 1449 -1848 3 gnd
rlabel metal1 1545 -1848 1545 -1848 7 vdd
rlabel metal1 1319 -1463 1319 -1463 5 vdd
rlabel metal1 1304 -1706 1304 -1706 1 gnd
rlabel metal1 1337 -1706 1337 -1706 1 gnd
rlabel metal1 1368 -1600 1368 -1600 5 vdd
rlabel metal1 1368 -1696 1368 -1696 1 gnd
rlabel metal1 1170 -1599 1170 -1599 5 vdd
rlabel metal1 1155 -1842 1155 -1842 1 gnd
rlabel metal1 1188 -1842 1188 -1842 1 gnd
rlabel metal1 1219 -1736 1219 -1736 5 vdd
rlabel metal1 1219 -1832 1219 -1832 1 gnd
rlabel metal1 1159 -1299 1159 -1299 5 vdd
rlabel metal1 1144 -1542 1144 -1542 1 gnd
rlabel metal1 1177 -1542 1177 -1542 1 gnd
rlabel metal1 1208 -1436 1208 -1436 5 vdd
rlabel metal1 1208 -1532 1208 -1532 1 gnd
rlabel metal1 1417 -2561 1417 -2561 1 gnd
rlabel metal1 1417 -2465 1417 -2465 5 vdd
rlabel metal1 1386 -2571 1386 -2571 1 gnd
rlabel metal1 1353 -2571 1353 -2571 1 gnd
rlabel metal1 1368 -2328 1368 -2328 5 vdd
rlabel metal1 1424 -2950 1424 -2950 1 gnd
rlabel metal1 1424 -2854 1424 -2854 5 vdd
rlabel metal1 1393 -2960 1393 -2960 1 gnd
rlabel metal1 1360 -2960 1360 -2960 1 gnd
rlabel metal1 1375 -2717 1375 -2717 5 vdd
rlabel metal1 1716 -3106 1716 -3106 1 gnd
rlabel metal1 1716 -3010 1716 -3010 5 vdd
rlabel metal1 1685 -3116 1685 -3116 1 gnd
rlabel metal1 1652 -3116 1652 -3116 1 gnd
rlabel metal1 1667 -2873 1667 -2873 5 vdd
rlabel metal1 2152 -2585 2152 -2585 1 gnd
rlabel metal1 2152 -2489 2152 -2489 5 vdd
rlabel metal1 2121 -2595 2121 -2595 1 gnd
rlabel metal1 2088 -2595 2088 -2595 1 gnd
rlabel metal1 2103 -2352 2103 -2352 5 vdd
rlabel metal1 762 -3055 762 -3055 1 gnd
rlabel metal1 762 -2959 762 -2959 5 vdd
rlabel metal1 719 -3086 719 -3086 1 gnd
rlabel metal1 727 -2889 727 -2889 5 vdd
rlabel metal1 700 -2889 700 -2889 5 vdd
rlabel metal1 766 -2784 766 -2784 1 gnd
rlabel metal1 766 -2688 766 -2688 5 vdd
rlabel metal1 723 -2815 723 -2815 1 gnd
rlabel metal1 731 -2618 731 -2618 5 vdd
rlabel metal1 704 -2618 704 -2618 5 vdd
rlabel metal1 765 -2501 765 -2501 1 gnd
rlabel metal1 765 -2405 765 -2405 5 vdd
rlabel metal1 722 -2532 722 -2532 1 gnd
rlabel metal1 730 -2335 730 -2335 5 vdd
rlabel metal1 703 -2335 703 -2335 5 vdd
rlabel metal1 750 -3304 750 -3304 1 gnd
rlabel metal1 750 -3208 750 -3208 5 vdd
rlabel metal1 715 -3138 715 -3138 5 vdd
rlabel metal1 688 -3138 688 -3138 5 vdd
rlabel metal1 707 -3335 707 -3335 1 gnd
rlabel metal1 1101 -2836 1101 -2836 1 gnd
rlabel metal1 1101 -2740 1101 -2740 5 vdd
rlabel metal1 1058 -2867 1058 -2867 1 gnd
rlabel metal1 1066 -2670 1066 -2670 5 vdd
rlabel metal1 1039 -2670 1039 -2670 5 vdd
rlabel metal1 1100 -2553 1100 -2553 1 gnd
rlabel metal1 1100 -2457 1100 -2457 5 vdd
rlabel metal1 1057 -2584 1057 -2584 1 gnd
rlabel metal1 1065 -2387 1065 -2387 5 vdd
rlabel metal1 1038 -2387 1038 -2387 5 vdd
rlabel metal1 767 -3571 767 -3571 1 gnd
rlabel metal1 767 -3475 767 -3475 5 vdd
rlabel metal1 724 -3602 724 -3602 1 gnd
rlabel metal1 732 -3405 732 -3405 5 vdd
rlabel metal1 705 -3405 705 -3405 5 vdd
rlabel metal1 755 -3820 755 -3820 1 gnd
rlabel metal1 755 -3724 755 -3724 5 vdd
rlabel metal1 720 -3654 720 -3654 5 vdd
rlabel metal1 693 -3654 693 -3654 5 vdd
rlabel metal1 712 -3851 712 -3851 1 gnd
rlabel metal1 1431 -3238 1431 -3238 1 gnd
rlabel metal1 1431 -3142 1431 -3142 5 vdd
rlabel metal1 1388 -3269 1388 -3269 1 gnd
rlabel metal1 1396 -3072 1396 -3072 5 vdd
rlabel metal1 1369 -3072 1369 -3072 5 vdd
rlabel metal1 1091 -3370 1091 -3370 1 gnd
rlabel metal1 1091 -3274 1091 -3274 5 vdd
rlabel metal1 1056 -3204 1056 -3204 5 vdd
rlabel metal1 1029 -3204 1029 -3204 5 vdd
rlabel metal1 1048 -3401 1048 -3401 1 gnd
rlabel metal1 -475 -89 -475 -89 1 clk
rlabel metal1 -253 98 -253 98 5 vdd
rlabel metal1 -254 -4 -254 -4 1 gnd
rlabel metal1 -221 98 -221 98 5 vdd
rlabel metal1 -222 -4 -222 -4 1 gnd
rlabel metal1 -298 90 -298 90 5 vdd
rlabel metal1 -298 -75 -298 -75 1 gnd
rlabel metal1 -350 90 -350 90 5 vdd
rlabel metal1 -350 -75 -350 -75 1 gnd
rlabel metal1 -402 -75 -402 -75 1 gnd
rlabel metal1 -402 90 -402 90 5 vdd
rlabel metal1 -454 -75 -454 -75 1 gnd
rlabel metal1 -454 90 -454 90 5 vdd
rlabel metal1 -442 -484 -442 -484 1 clk
rlabel metal1 -220 -297 -220 -297 5 vdd
rlabel metal1 -221 -399 -221 -399 1 gnd
rlabel metal1 -188 -297 -188 -297 5 vdd
rlabel metal1 -189 -399 -189 -399 1 gnd
rlabel metal1 -265 -305 -265 -305 5 vdd
rlabel metal1 -265 -470 -265 -470 1 gnd
rlabel metal1 -317 -305 -317 -305 5 vdd
rlabel metal1 -317 -470 -317 -470 1 gnd
rlabel metal1 -369 -470 -369 -470 1 gnd
rlabel metal1 -369 -305 -369 -305 5 vdd
rlabel metal1 -421 -470 -421 -470 1 gnd
rlabel metal1 -421 -305 -421 -305 5 vdd
rlabel metal1 -551 -863 -551 -863 1 clk
rlabel metal1 -329 -676 -329 -676 5 vdd
rlabel metal1 -330 -778 -330 -778 1 gnd
rlabel metal1 -297 -676 -297 -676 5 vdd
rlabel metal1 -298 -778 -298 -778 1 gnd
rlabel metal1 -374 -684 -374 -684 5 vdd
rlabel metal1 -374 -849 -374 -849 1 gnd
rlabel metal1 -426 -684 -426 -684 5 vdd
rlabel metal1 -426 -849 -426 -849 1 gnd
rlabel metal1 -478 -849 -478 -849 1 gnd
rlabel metal1 -478 -684 -478 -684 5 vdd
rlabel metal1 -530 -849 -530 -849 1 gnd
rlabel metal1 -530 -684 -530 -684 5 vdd
rlabel metal1 -454 -1037 -454 -1037 5 vdd
rlabel metal1 -454 -1202 -454 -1202 1 gnd
rlabel metal1 -402 -1037 -402 -1037 5 vdd
rlabel metal1 -402 -1202 -402 -1202 1 gnd
rlabel metal1 -350 -1202 -350 -1202 1 gnd
rlabel metal1 -350 -1037 -350 -1037 5 vdd
rlabel metal1 -298 -1202 -298 -1202 1 gnd
rlabel metal1 -298 -1037 -298 -1037 5 vdd
rlabel metal1 -222 -1131 -222 -1131 1 gnd
rlabel metal1 -221 -1029 -221 -1029 5 vdd
rlabel metal1 -254 -1131 -254 -1131 1 gnd
rlabel metal1 -253 -1029 -253 -1029 5 vdd
rlabel metal1 -475 -1216 -475 -1216 1 clk
rlabel metal1 -463 -1365 -463 -1365 5 vdd
rlabel metal1 -463 -1530 -463 -1530 1 gnd
rlabel metal1 -411 -1365 -411 -1365 5 vdd
rlabel metal1 -411 -1530 -411 -1530 1 gnd
rlabel metal1 -359 -1530 -359 -1530 1 gnd
rlabel metal1 -359 -1365 -359 -1365 5 vdd
rlabel metal1 -307 -1530 -307 -1530 1 gnd
rlabel metal1 -307 -1365 -307 -1365 5 vdd
rlabel metal1 -231 -1459 -231 -1459 1 gnd
rlabel metal1 -230 -1357 -230 -1357 5 vdd
rlabel metal1 -263 -1459 -263 -1459 1 gnd
rlabel metal1 -262 -1357 -262 -1357 5 vdd
rlabel metal1 -484 -1544 -484 -1544 1 clk
rlabel metal1 -500 -1922 -500 -1922 1 clk
rlabel metal1 -278 -1735 -278 -1735 5 vdd
rlabel metal1 -279 -1837 -279 -1837 1 gnd
rlabel metal1 -246 -1735 -246 -1735 5 vdd
rlabel metal1 -247 -1837 -247 -1837 1 gnd
rlabel metal1 -323 -1743 -323 -1743 5 vdd
rlabel metal1 -323 -1908 -323 -1908 1 gnd
rlabel metal1 -375 -1743 -375 -1743 5 vdd
rlabel metal1 -375 -1908 -375 -1908 1 gnd
rlabel metal1 -427 -1908 -427 -1908 1 gnd
rlabel metal1 -427 -1743 -427 -1743 5 vdd
rlabel metal1 -479 -1908 -479 -1908 1 gnd
rlabel metal1 -479 -1743 -479 -1743 5 vdd
rlabel metal1 -484 -2292 -484 -2292 1 clk
rlabel metal1 -262 -2105 -262 -2105 5 vdd
rlabel metal1 -263 -2207 -263 -2207 1 gnd
rlabel metal1 -230 -2105 -230 -2105 5 vdd
rlabel metal1 -231 -2207 -231 -2207 1 gnd
rlabel metal1 -307 -2113 -307 -2113 5 vdd
rlabel metal1 -307 -2278 -307 -2278 1 gnd
rlabel metal1 -359 -2113 -359 -2113 5 vdd
rlabel metal1 -359 -2278 -359 -2278 1 gnd
rlabel metal1 -411 -2278 -411 -2278 1 gnd
rlabel metal1 -411 -2113 -411 -2113 5 vdd
rlabel metal1 -463 -2278 -463 -2278 1 gnd
rlabel metal1 -463 -2113 -463 -2113 5 vdd
rlabel metal1 -475 -2721 -475 -2721 1 clk
rlabel metal1 -253 -2534 -253 -2534 5 vdd
rlabel metal1 -254 -2636 -254 -2636 1 gnd
rlabel metal1 -221 -2534 -221 -2534 5 vdd
rlabel metal1 -222 -2636 -222 -2636 1 gnd
rlabel metal1 -298 -2542 -298 -2542 5 vdd
rlabel metal1 -298 -2707 -298 -2707 1 gnd
rlabel metal1 -350 -2542 -350 -2542 5 vdd
rlabel metal1 -350 -2707 -350 -2707 1 gnd
rlabel metal1 -402 -2707 -402 -2707 1 gnd
rlabel metal1 -402 -2542 -402 -2542 5 vdd
rlabel metal1 -454 -2707 -454 -2707 1 gnd
rlabel metal1 -454 -2542 -454 -2542 5 vdd
rlabel metal1 1156 37 1156 37 1 clk
rlabel metal1 1378 224 1378 224 5 vdd
rlabel metal1 1377 122 1377 122 1 gnd
rlabel metal1 1410 224 1410 224 5 vdd
rlabel metal1 1409 122 1409 122 1 gnd
rlabel metal1 1333 216 1333 216 5 vdd
rlabel metal1 1333 51 1333 51 1 gnd
rlabel metal1 1281 216 1281 216 5 vdd
rlabel metal1 1281 51 1281 51 1 gnd
rlabel metal1 1229 51 1229 51 1 gnd
rlabel metal1 1229 216 1229 216 5 vdd
rlabel metal1 1177 51 1177 51 1 gnd
rlabel metal1 1177 216 1177 216 5 vdd
rlabel metal1 1434 -426 1434 -426 1 clk
rlabel metal1 1656 -239 1656 -239 5 vdd
rlabel metal1 1655 -341 1655 -341 1 gnd
rlabel metal1 1688 -239 1688 -239 5 vdd
rlabel metal1 1687 -341 1687 -341 1 gnd
rlabel metal1 1611 -247 1611 -247 5 vdd
rlabel metal1 1611 -412 1611 -412 1 gnd
rlabel metal1 1559 -247 1559 -247 5 vdd
rlabel metal1 1559 -412 1559 -412 1 gnd
rlabel metal1 1507 -412 1507 -412 1 gnd
rlabel metal1 1507 -247 1507 -247 5 vdd
rlabel metal1 1455 -412 1455 -412 1 gnd
rlabel metal1 1455 -247 1455 -247 5 vdd
rlabel metal1 1745 -981 1745 -981 1 clk
rlabel metal1 1967 -794 1967 -794 5 vdd
rlabel metal1 1966 -896 1966 -896 1 gnd
rlabel metal1 1999 -794 1999 -794 5 vdd
rlabel metal1 1998 -896 1998 -896 1 gnd
rlabel metal1 1922 -802 1922 -802 5 vdd
rlabel metal1 1922 -967 1922 -967 1 gnd
rlabel metal1 1870 -802 1870 -802 5 vdd
rlabel metal1 1870 -967 1870 -967 1 gnd
rlabel metal1 1818 -967 1818 -967 1 gnd
rlabel metal1 1818 -802 1818 -802 5 vdd
rlabel metal1 1766 -967 1766 -967 1 gnd
rlabel metal1 1766 -802 1766 -802 5 vdd
rlabel metal1 1896 -1931 1896 -1931 1 clk
rlabel metal1 2118 -1744 2118 -1744 5 vdd
rlabel metal1 2117 -1846 2117 -1846 1 gnd
rlabel metal1 2150 -1744 2150 -1744 5 vdd
rlabel metal1 2149 -1846 2149 -1846 1 gnd
rlabel metal1 2073 -1752 2073 -1752 5 vdd
rlabel metal1 2073 -1917 2073 -1917 1 gnd
rlabel metal1 2021 -1752 2021 -1752 5 vdd
rlabel metal1 2021 -1917 2021 -1917 1 gnd
rlabel metal1 1969 -1917 1969 -1917 1 gnd
rlabel metal1 1969 -1752 1969 -1752 5 vdd
rlabel metal1 1917 -1917 1917 -1917 1 gnd
rlabel metal1 1917 -1752 1917 -1752 5 vdd
rlabel metal1 2426 -2612 2426 -2612 1 clk
rlabel metal1 2648 -2425 2648 -2425 5 vdd
rlabel metal1 2647 -2527 2647 -2527 1 gnd
rlabel metal1 2680 -2425 2680 -2425 5 vdd
rlabel metal1 2679 -2527 2679 -2527 1 gnd
rlabel metal1 2603 -2433 2603 -2433 5 vdd
rlabel metal1 2603 -2598 2603 -2598 1 gnd
rlabel metal1 2551 -2433 2551 -2433 5 vdd
rlabel metal1 2551 -2598 2551 -2598 1 gnd
rlabel metal1 2499 -2598 2499 -2598 1 gnd
rlabel metal1 2499 -2433 2499 -2433 5 vdd
rlabel metal1 2447 -2598 2447 -2598 1 gnd
rlabel metal1 2447 -2433 2447 -2433 5 vdd
rlabel metal1 -481 8 -481 8 1 A0
rlabel metal1 -210 32 -210 32 1 A_D0
rlabel metal1 -14 -174 -14 -174 1 A_D0
rlabel metal1 -448 -394 -448 -394 1 B0
rlabel metal1 -176 -362 -176 -362 1 B_D0
rlabel metal1 -13 -222 -13 -222 1 B_D0
rlabel metal1 -558 -764 -558 -764 3 A1
rlabel metal1 -285 -743 -285 -743 1 A_D1
rlabel metal1 -481 -1137 -481 -1137 1 B1
rlabel metal1 -209 -1095 -209 -1095 1 B_D1
rlabel metal1 -63 -810 -63 -810 1 A_D1
rlabel metal1 -58 -858 -58 -858 1 B_D1
rlabel metal1 -219 -1423 -219 -1423 1 A_D2
rlabel metal1 -490 -1442 -490 -1442 1 A2
rlabel metal1 -506 -1820 -506 -1820 1 B2
rlabel metal1 -234 -1801 -234 -1801 1 B_D2
rlabel metal1 -52 -1470 -52 -1470 1 A_D2
rlabel metal1 -54 -1518 -54 -1518 1 B_D2
rlabel metal1 -489 -2214 -489 -2214 1 A3
rlabel metal1 -220 -2171 -220 -2171 1 A_D3
rlabel metal1 -209 -2600 -209 -2600 1 B_D3
rlabel metal1 -481 -2630 -481 -2630 1 B3
rlabel metal1 -58 -2345 -58 -2345 1 A_D3
rlabel metal1 -54 -2391 -54 -2391 1 B_D3
rlabel metal1 665 -25 665 -25 1 S_D0
rlabel metal1 1150 141 1150 141 1 S_D0
rlabel metal1 1421 158 1421 158 1 S0
rlabel metal1 1156 -411 1156 -411 1 S_D1
rlabel metal1 1427 -344 1427 -344 1 S_D1
rlabel metal1 1702 -304 1702 -304 1 S1
rlabel metal1 1493 -857 1493 -857 1 S_D2
rlabel metal1 1739 -891 1739 -891 1 S_D2
rlabel metal1 2010 -861 2010 -861 1 S2
rlabel metal1 1607 -1821 1607 -1821 1 S_D3
rlabel metal1 1891 -1858 1891 -1858 1 S_D3
rlabel metal1 2162 -1810 2162 -1810 1 S3
rlabel metal1 2184 -2551 2184 -2551 1 c_d4
rlabel metal1 2421 -2532 2421 -2532 1 c_d4
rlabel metal1 2693 -2491 2693 -2491 7 c4
<< end >>
